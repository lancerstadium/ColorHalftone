/**
 * Module       : LUTTable
 * Input        : x[7:0] - Signed/Unsigned 8-bit interger
 * Output       : y[7:0] - Unsigned/Signed 8-bit interger
 * Description  : LUT Table for read and write.
 * Author       : lancerstadium
 * Date         : Sat Mar  1 00:00:00 CST 2025
 * License      : MIT
 */

module LUTTable_x4_4b_i8_s1_D_H6 (
    // 系统接口
    input  logic         clk,      // 全局时钟
    input  logic         rst_n,    // 异步复位
    // 批量读取控制
    input  logic         burst_start,  // 脉冲启动批量读取
    output logic         burst_done,   // 批量读取完成标志
    input  logic [13:0] base_addr,  // 展平后基地址
    // 数据输出
    output logic signed [7:0] data [0:15]  // 并行输出
);

    (* rom_style = "block" *) 
    logic signed [7:0] lut_mem [0:9215]
    // Original Shape: (576, 16), Total Entries: 9216
'{
    /* (0, 0) */	    8'shfb, 8'sh0b, 8'sh19, 8'she1, 8'sh11, 8'shf3, 8'she7, 8'shfe, 8'sh03, 8'shea, 8'sh07, 8'shfd, 8'sh0e, 8'shfd, 8'sh1a, 8'shfe
    /* (1, 0) */	    8'shfc, 8'sh0b, 8'sh18, 8'she2, 8'sh10, 8'shf4, 8'she7, 8'shfe, 8'sh03, 8'sheb, 8'sh07, 8'shfd, 8'sh0e, 8'shfd, 8'sh19, 8'shfe
    /* (2, 0) */	    8'shfc, 8'sh0a, 8'sh18, 8'she3, 8'sh10, 8'shf4, 8'she8, 8'shfe, 8'sh03, 8'shec, 8'sh07, 8'shfd, 8'sh0e, 8'shfe, 8'sh18, 8'shfe
    /* (3, 0) */	    8'shfc, 8'sh0a, 8'sh17, 8'she4, 8'sh0f, 8'shf5, 8'she9, 8'shfe, 8'sh03, 8'shec, 8'sh07, 8'shfe, 8'sh0d, 8'shfe, 8'sh17, 8'shff
    /* (4, 0) */	    8'shfc, 8'sh09, 8'sh16, 8'she5, 8'sh0f, 8'shf5, 8'shea, 8'shfe, 8'sh03, 8'shed, 8'sh07, 8'shfe, 8'sh0d, 8'shfe, 8'sh17, 8'shff
    /* (5, 0) */	    8'shfc, 8'sh09, 8'sh15, 8'she5, 8'sh0e, 8'shf5, 8'sheb, 8'shfe, 8'sh03, 8'shee, 8'sh06, 8'shfe, 8'sh0c, 8'shfe, 8'sh16, 8'shff
    /* (6, 0) */	    8'shfc, 8'sh09, 8'sh14, 8'she6, 8'sh0e, 8'shf6, 8'sheb, 8'shfe, 8'sh03, 8'shee, 8'sh06, 8'shfe, 8'sh0c, 8'shfe, 8'sh15, 8'shff
    /* (7, 0) */	    8'shfc, 8'sh08, 8'sh14, 8'she7, 8'sh0d, 8'shf6, 8'shec, 8'shfe, 8'sh02, 8'shef, 8'sh06, 8'shfe, 8'sh0b, 8'shfe, 8'sh14, 8'shff
    /* (8, 0) */	    8'shfd, 8'sh08, 8'sh13, 8'she8, 8'sh0d, 8'shf7, 8'shed, 8'shfe, 8'sh02, 8'shf0, 8'sh06, 8'shfe, 8'sh0b, 8'shfe, 8'sh13, 8'shff
    /* (9, 0) */	    8'shfd, 8'sh08, 8'sh12, 8'she9, 8'sh0c, 8'shf7, 8'shee, 8'shfe, 8'sh02, 8'shf0, 8'sh05, 8'shfe, 8'sh0a, 8'shfe, 8'sh13, 8'shff
    /* (10, 0) */	    8'shfd, 8'sh07, 8'sh11, 8'shea, 8'sh0c, 8'shf7, 8'shef, 8'shfe, 8'sh02, 8'shf1, 8'sh05, 8'shfe, 8'sh0a, 8'shfe, 8'sh12, 8'shff
    /* (11, 0) */	    8'shfd, 8'sh07, 8'sh11, 8'sheb, 8'sh0b, 8'shf8, 8'shef, 8'shfe, 8'sh02, 8'shf2, 8'sh05, 8'shfe, 8'sh09, 8'shfe, 8'sh11, 8'shff
    /* (12, 0) */	    8'shfd, 8'sh07, 8'sh10, 8'shec, 8'sh0b, 8'shf8, 8'shf0, 8'shfe, 8'sh02, 8'shf2, 8'sh05, 8'shfe, 8'sh09, 8'shfe, 8'sh10, 8'shff
    /* (13, 0) */	    8'shfd, 8'sh06, 8'sh0f, 8'shed, 8'sh0a, 8'shf9, 8'shf1, 8'shff, 8'sh02, 8'shf3, 8'sh04, 8'shfe, 8'sh09, 8'shfe, 8'sh0f, 8'shff
    /* (14, 0) */	    8'shfd, 8'sh06, 8'sh0e, 8'shee, 8'sh0a, 8'shf9, 8'shf2, 8'shff, 8'sh02, 8'shf4, 8'sh04, 8'shfe, 8'sh08, 8'shff, 8'sh0f, 8'shff
    /* (15, 0) */	    8'shfe, 8'sh06, 8'sh0d, 8'shef, 8'sh09, 8'shf9, 8'shf3, 8'shff, 8'sh02, 8'shf4, 8'sh04, 8'shff, 8'sh08, 8'shff, 8'sh0e, 8'shff
    /* (16, 0) */	    8'shfe, 8'sh05, 8'sh0d, 8'shf0, 8'sh08, 8'shfa, 8'shf3, 8'shff, 8'sh02, 8'shf5, 8'sh04, 8'shff, 8'sh07, 8'shff, 8'sh0d, 8'shff
    /* (17, 0) */	    8'shfe, 8'sh05, 8'sh0c, 8'shf1, 8'sh08, 8'shfa, 8'shf4, 8'shff, 8'sh01, 8'shf6, 8'sh04, 8'shff, 8'sh07, 8'shff, 8'sh0c, 8'shff
    /* (18, 0) */	    8'shfe, 8'sh05, 8'sh0b, 8'shf2, 8'sh07, 8'shfa, 8'shf5, 8'shff, 8'sh01, 8'shf6, 8'sh03, 8'shff, 8'sh06, 8'shff, 8'sh0b, 8'shff
    /* (19, 0) */	    8'shfe, 8'sh04, 8'sh0a, 8'shf3, 8'sh07, 8'shfb, 8'shf6, 8'shff, 8'sh01, 8'shf7, 8'sh03, 8'shff, 8'sh06, 8'shff, 8'sh0b, 8'shff
    /* (20, 0) */	    8'shfe, 8'sh04, 8'sh09, 8'shf4, 8'sh06, 8'shfb, 8'shf6, 8'shff, 8'sh01, 8'shf8, 8'sh03, 8'shff, 8'sh05, 8'shff, 8'sh0a, 8'shff
    /* (21, 0) */	    8'shfe, 8'sh04, 8'sh09, 8'shf5, 8'sh06, 8'shfc, 8'shf7, 8'shff, 8'sh01, 8'shf9, 8'sh03, 8'shff, 8'sh05, 8'shff, 8'sh09, 8'shff
    /* (22, 0) */	    8'shff, 8'sh03, 8'sh08, 8'shf6, 8'sh05, 8'shfc, 8'shf8, 8'shff, 8'sh01, 8'shf9, 8'sh02, 8'shff, 8'sh05, 8'shff, 8'sh08, 8'shff
    /* (23, 0) */	    8'shff, 8'sh03, 8'sh07, 8'shf7, 8'sh05, 8'shfc, 8'shf9, 8'shff, 8'sh01, 8'shfa, 8'sh02, 8'shff, 8'sh04, 8'shff, 8'sh07, 8'sh00
    /* (24, 0) */	    8'shff, 8'sh03, 8'sh06, 8'shf8, 8'sh04, 8'shfd, 8'shfa, 8'shff, 8'sh01, 8'shfb, 8'sh02, 8'shff, 8'sh04, 8'shff, 8'sh06, 8'sh00
    /* (25, 0) */	    8'shff, 8'sh02, 8'sh06, 8'shf9, 8'sh04, 8'shfd, 8'shfa, 8'shff, 8'sh01, 8'shfb, 8'sh02, 8'shff, 8'sh03, 8'shff, 8'sh06, 8'sh00
    /* (26, 0) */	    8'shff, 8'sh02, 8'sh05, 8'shfa, 8'sh03, 8'shfe, 8'shfb, 8'sh00, 8'sh01, 8'shfc, 8'sh01, 8'shff, 8'sh03, 8'sh00, 8'sh05, 8'sh00
    /* (27, 0) */	    8'shff, 8'sh02, 8'sh04, 8'shfb, 8'sh03, 8'shfe, 8'shfc, 8'sh00, 8'sh00, 8'shfd, 8'sh01, 8'sh00, 8'sh02, 8'sh00, 8'sh04, 8'sh00
    /* (28, 0) */	    8'shff, 8'sh01, 8'sh03, 8'shfc, 8'sh02, 8'shfe, 8'shfd, 8'sh00, 8'sh00, 8'shfd, 8'sh01, 8'sh00, 8'sh02, 8'sh00, 8'sh03, 8'sh00
    /* (29, 0) */	    8'sh00, 8'sh01, 8'sh02, 8'shfd, 8'sh02, 8'shff, 8'shfe, 8'sh00, 8'sh00, 8'shfe, 8'sh01, 8'sh00, 8'sh01, 8'sh00, 8'sh02, 8'sh00
    /* (30, 0) */	    8'sh00, 8'sh01, 8'sh02, 8'shfe, 8'sh01, 8'shff, 8'shfe, 8'sh00, 8'sh00, 8'shff, 8'sh00, 8'sh00, 8'sh01, 8'sh00, 8'sh02, 8'sh00
    /* (31, 0) */	    8'sh00, 8'sh00, 8'sh01, 8'shff, 8'sh01, 8'sh00, 8'shff, 8'sh00, 8'sh00, 8'shff, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh01, 8'sh00
    /* (32, 0) */	    8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00
    /* (33, 0) */	    8'sh00, 8'sh00, 8'shff, 8'sh01, 8'shff, 8'sh00, 8'sh01, 8'sh00, 8'sh00, 8'sh01, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'shff, 8'sh00
    /* (34, 0) */	    8'sh00, 8'shff, 8'shfe, 8'sh02, 8'shff, 8'sh01, 8'sh02, 8'sh00, 8'sh00, 8'sh01, 8'sh00, 8'sh00, 8'shff, 8'sh00, 8'shfe, 8'sh00
    /* (35, 0) */	    8'sh00, 8'shff, 8'shfe, 8'sh03, 8'shfe, 8'sh01, 8'sh02, 8'sh00, 8'sh00, 8'sh02, 8'shff, 8'sh00, 8'shff, 8'sh00, 8'shfe, 8'sh00
    /* (36, 0) */	    8'sh01, 8'shff, 8'shfd, 8'sh04, 8'shfe, 8'sh02, 8'sh03, 8'sh00, 8'sh00, 8'sh03, 8'shff, 8'sh00, 8'shfe, 8'sh00, 8'shfd, 8'sh00
    /* (37, 0) */	    8'sh01, 8'shfe, 8'shfc, 8'sh05, 8'shfd, 8'sh02, 8'sh04, 8'sh00, 8'sh00, 8'sh03, 8'shff, 8'sh00, 8'shfe, 8'sh00, 8'shfc, 8'sh00
    /* (38, 0) */	    8'sh01, 8'shfe, 8'shfb, 8'sh06, 8'shfd, 8'sh02, 8'sh05, 8'sh00, 8'shff, 8'sh04, 8'shff, 8'sh01, 8'shfd, 8'sh00, 8'shfb, 8'sh00
    /* (39, 0) */	    8'sh01, 8'shfe, 8'shfa, 8'sh07, 8'shfc, 8'sh03, 8'sh06, 8'sh01, 8'shff, 8'sh05, 8'shfe, 8'sh01, 8'shfd, 8'sh01, 8'shfa, 8'sh00
    /* (40, 0) */	    8'sh01, 8'shfd, 8'shfa, 8'sh08, 8'shfc, 8'sh03, 8'sh06, 8'sh01, 8'shff, 8'sh05, 8'shfe, 8'sh01, 8'shfc, 8'sh01, 8'shfa, 8'sh00
    /* (41, 0) */	    8'sh01, 8'shfd, 8'shf9, 8'sh09, 8'shfb, 8'sh04, 8'sh07, 8'sh01, 8'shff, 8'sh06, 8'shfe, 8'sh01, 8'shfc, 8'sh01, 8'shf9, 8'sh00
    /* (42, 0) */	    8'sh01, 8'shfd, 8'shf8, 8'sh0a, 8'shfb, 8'sh04, 8'sh08, 8'sh01, 8'shff, 8'sh07, 8'shfe, 8'sh01, 8'shfb, 8'sh01, 8'shf8, 8'sh01
    /* (43, 0) */	    8'sh02, 8'shfc, 8'shf7, 8'sh0b, 8'shfa, 8'sh04, 8'sh09, 8'sh01, 8'shff, 8'sh07, 8'shfd, 8'sh01, 8'shfb, 8'sh01, 8'shf7, 8'sh01
    /* (44, 0) */	    8'sh02, 8'shfc, 8'shf7, 8'sh0c, 8'shfa, 8'sh05, 8'sh0a, 8'sh01, 8'shff, 8'sh08, 8'shfd, 8'sh01, 8'shfb, 8'sh01, 8'shf6, 8'sh01
    /* (45, 0) */	    8'sh02, 8'shfc, 8'shf6, 8'sh0d, 8'shf9, 8'sh05, 8'sh0a, 8'sh01, 8'shff, 8'sh09, 8'shfd, 8'sh01, 8'shfa, 8'sh01, 8'shf5, 8'sh01
    /* (46, 0) */	    8'sh02, 8'shfb, 8'shf5, 8'sh0e, 8'shf9, 8'sh06, 8'sh0b, 8'sh01, 8'shff, 8'sh0a, 8'shfd, 8'sh01, 8'shfa, 8'sh01, 8'shf5, 8'sh01
    /* (47, 0) */	    8'sh02, 8'shfb, 8'shf4, 8'sh0f, 8'shf8, 8'sh06, 8'sh0c, 8'sh01, 8'shff, 8'sh0a, 8'shfc, 8'sh01, 8'shf9, 8'sh01, 8'shf4, 8'sh01
    /* (48, 0) */	    8'sh02, 8'shfb, 8'shf3, 8'sh10, 8'shf8, 8'sh06, 8'sh0d, 8'sh01, 8'shfe, 8'sh0b, 8'shfc, 8'sh01, 8'shf9, 8'sh01, 8'shf3, 8'sh01
    /* (49, 0) */	    8'sh02, 8'shfa, 8'shf3, 8'sh11, 8'shf7, 8'sh07, 8'sh0d, 8'sh01, 8'shfe, 8'sh0c, 8'shfc, 8'sh01, 8'shf8, 8'sh01, 8'shf2, 8'sh01
    /* (50, 0) */	    8'sh03, 8'shfa, 8'shf2, 8'sh12, 8'shf6, 8'sh07, 8'sh0e, 8'sh01, 8'shfe, 8'sh0c, 8'shfc, 8'sh02, 8'shf8, 8'sh01, 8'shf1, 8'sh01
    /* (51, 0) */	    8'sh03, 8'shfa, 8'shf1, 8'sh13, 8'shf6, 8'sh07, 8'sh0f, 8'sh01, 8'shfe, 8'sh0d, 8'shfc, 8'sh02, 8'shf7, 8'sh02, 8'shf1, 8'sh01
    /* (52, 0) */	    8'sh03, 8'shf9, 8'shf0, 8'sh14, 8'shf5, 8'sh08, 8'sh10, 8'sh02, 8'shfe, 8'sh0e, 8'shfb, 8'sh02, 8'shf7, 8'sh02, 8'shf0, 8'sh01
    /* (53, 0) */	    8'sh03, 8'shf9, 8'shef, 8'sh15, 8'shf5, 8'sh08, 8'sh11, 8'sh02, 8'shfe, 8'sh0e, 8'shfb, 8'sh02, 8'shf7, 8'sh02, 8'shef, 8'sh01
    /* (54, 0) */	    8'sh03, 8'shf9, 8'shef, 8'sh16, 8'shf4, 8'sh09, 8'sh11, 8'sh02, 8'shfe, 8'sh0f, 8'shfb, 8'sh02, 8'shf6, 8'sh02, 8'shee, 8'sh01
    /* (55, 0) */	    8'sh03, 8'shf8, 8'shee, 8'sh17, 8'shf4, 8'sh09, 8'sh12, 8'sh02, 8'shfe, 8'sh10, 8'shfb, 8'sh02, 8'shf6, 8'sh02, 8'shed, 8'sh01
    /* (56, 0) */	    8'sh03, 8'shf8, 8'shed, 8'sh18, 8'shf3, 8'sh09, 8'sh13, 8'sh02, 8'shfe, 8'sh10, 8'shfa, 8'sh02, 8'shf5, 8'sh02, 8'shed, 8'sh01
    /* (57, 0) */	    8'sh04, 8'shf8, 8'shec, 8'sh19, 8'shf3, 8'sh0a, 8'sh14, 8'sh02, 8'shfe, 8'sh11, 8'shfa, 8'sh02, 8'shf5, 8'sh02, 8'shec, 8'sh01
    /* (58, 0) */	    8'sh04, 8'shf7, 8'shec, 8'sh1a, 8'shf2, 8'sh0a, 8'sh15, 8'sh02, 8'shfd, 8'sh12, 8'shfa, 8'sh02, 8'shf4, 8'sh02, 8'sheb, 8'sh01
    /* (59, 0) */	    8'sh04, 8'shf7, 8'sheb, 8'sh1b, 8'shf2, 8'sh0b, 8'sh15, 8'sh02, 8'shfd, 8'sh12, 8'shfa, 8'sh02, 8'shf4, 8'sh02, 8'shea, 8'sh01
    /* (60, 0) */	    8'sh04, 8'shf7, 8'shea, 8'sh1b, 8'shf1, 8'sh0b, 8'sh16, 8'sh02, 8'shfd, 8'sh13, 8'shf9, 8'sh02, 8'shf3, 8'sh02, 8'she9, 8'sh01
    /* (61, 0) */	    8'sh04, 8'shf6, 8'she9, 8'sh1c, 8'shf1, 8'sh0b, 8'sh17, 8'sh02, 8'shfd, 8'sh14, 8'shf9, 8'sh02, 8'shf3, 8'sh02, 8'she9, 8'sh01
    /* (62, 0) */	    8'sh04, 8'shf6, 8'she8, 8'sh1d, 8'shf0, 8'sh0c, 8'sh18, 8'sh02, 8'shfd, 8'sh14, 8'shf9, 8'sh03, 8'shf2, 8'sh02, 8'she8, 8'sh02
    /* (63, 0) */	    8'sh04, 8'shf5, 8'she8, 8'sh1e, 8'shf0, 8'sh0c, 8'sh19, 8'sh02, 8'shfd, 8'sh15, 8'shf9, 8'sh03, 8'shf2, 8'sh03, 8'she7, 8'sh02
    /* (64, 0) */	    8'sh09, 8'shf4, 8'shdf, 8'sh12, 8'shf5, 8'sh43, 8'shed, 8'she9, 8'shf8, 8'sh08, 8'shff, 8'sh50, 8'shf2, 8'shf3, 8'shd0, 8'sh32
    /* (65, 0) */	    8'sh09, 8'shf4, 8'she1, 8'sh12, 8'shf5, 8'sh41, 8'shed, 8'shea, 8'shf8, 8'sh08, 8'shff, 8'sh4d, 8'shf2, 8'shf4, 8'shd1, 8'sh30
    /* (66, 0) */	    8'sh09, 8'shf5, 8'she2, 8'sh11, 8'shf5, 8'sh3f, 8'shee, 8'sheb, 8'shf8, 8'sh07, 8'shff, 8'sh4b, 8'shf3, 8'shf4, 8'shd3, 8'sh2e
    /* (67, 0) */	    8'sh08, 8'shf5, 8'she3, 8'sh11, 8'shf6, 8'sh3d, 8'shee, 8'sheb, 8'shf8, 8'sh07, 8'shff, 8'sh48, 8'shf3, 8'shf4, 8'shd4, 8'sh2d
    /* (68, 0) */	    8'sh08, 8'shf6, 8'she4, 8'sh10, 8'shf6, 8'sh3b, 8'shef, 8'shec, 8'shf9, 8'sh07, 8'shff, 8'sh46, 8'shf4, 8'shf5, 8'shd6, 8'sh2b
    /* (69, 0) */	    8'sh08, 8'shf6, 8'she5, 8'sh0f, 8'shf6, 8'sh39, 8'shf0, 8'shed, 8'shf9, 8'sh07, 8'shff, 8'sh43, 8'shf4, 8'shf5, 8'shd7, 8'sh2a
    /* (70, 0) */	    8'sh07, 8'shf6, 8'she6, 8'sh0f, 8'shf7, 8'sh36, 8'shf0, 8'shed, 8'shf9, 8'sh06, 8'shff, 8'sh41, 8'shf5, 8'shf6, 8'shd9, 8'sh28
    /* (71, 0) */	    8'sh07, 8'shf7, 8'she7, 8'sh0e, 8'shf7, 8'sh34, 8'shf1, 8'shee, 8'shf9, 8'sh06, 8'shff, 8'sh3e, 8'shf5, 8'shf6, 8'shda, 8'sh27
    /* (72, 0) */	    8'sh07, 8'shf7, 8'she8, 8'sh0e, 8'shf7, 8'sh32, 8'shf1, 8'shef, 8'shfa, 8'sh06, 8'shff, 8'sh3c, 8'shf6, 8'shf6, 8'shdc, 8'sh25
    /* (73, 0) */	    8'sh07, 8'shf7, 8'she9, 8'sh0d, 8'shf8, 8'sh30, 8'shf2, 8'shf0, 8'shfa, 8'sh06, 8'shff, 8'sh39, 8'shf6, 8'shf7, 8'shdd, 8'sh24
    /* (74, 0) */	    8'sh06, 8'shf8, 8'shea, 8'sh0d, 8'shf8, 8'sh2e, 8'shf3, 8'shf0, 8'shfa, 8'sh05, 8'shff, 8'sh37, 8'shf6, 8'shf7, 8'shdf, 8'sh22
    /* (75, 0) */	    8'sh06, 8'shf8, 8'sheb, 8'sh0c, 8'shf8, 8'sh2c, 8'shf3, 8'shf1, 8'shfa, 8'sh05, 8'sh00, 8'sh34, 8'shf7, 8'shf8, 8'she0, 8'sh21
    /* (76, 0) */	    8'sh06, 8'shf9, 8'shec, 8'sh0b, 8'shf9, 8'sh2a, 8'shf4, 8'shf2, 8'shfb, 8'sh05, 8'sh00, 8'sh32, 8'shf7, 8'shf8, 8'she2, 8'sh1f
    /* (77, 0) */	    8'sh05, 8'shf9, 8'shed, 8'sh0b, 8'shf9, 8'sh28, 8'shf4, 8'shf2, 8'shfb, 8'sh05, 8'sh00, 8'sh2f, 8'shf8, 8'shf8, 8'she3, 8'sh1d
    /* (78, 0) */	    8'sh05, 8'shf9, 8'shee, 8'sh0a, 8'shfa, 8'sh26, 8'shf5, 8'shf3, 8'shfb, 8'sh04, 8'sh00, 8'sh2d, 8'shf8, 8'shf9, 8'she5, 8'sh1c
    /* (79, 0) */	    8'sh05, 8'shfa, 8'shef, 8'sh0a, 8'shfa, 8'sh24, 8'shf6, 8'shf4, 8'shfb, 8'sh04, 8'sh00, 8'sh2a, 8'shf9, 8'shf9, 8'she6, 8'sh1a
    /* (80, 0) */	    8'sh05, 8'shfa, 8'shf0, 8'sh09, 8'shfa, 8'sh22, 8'shf6, 8'shf5, 8'shfc, 8'sh04, 8'sh00, 8'sh28, 8'shf9, 8'shfa, 8'she8, 8'sh19
    /* (81, 0) */	    8'sh04, 8'shfa, 8'shf1, 8'sh09, 8'shfb, 8'sh1f, 8'shf7, 8'shf5, 8'shfc, 8'sh04, 8'sh00, 8'sh25, 8'shf9, 8'shfa, 8'she9, 8'sh17
    /* (82, 0) */	    8'sh04, 8'shfb, 8'shf2, 8'sh08, 8'shfb, 8'sh1d, 8'shf7, 8'shf6, 8'shfc, 8'sh03, 8'sh00, 8'sh23, 8'shfa, 8'shfa, 8'sheb, 8'sh16
    /* (83, 0) */	    8'sh04, 8'shfb, 8'shf3, 8'sh07, 8'shfb, 8'sh1b, 8'shf8, 8'shf7, 8'shfd, 8'sh03, 8'sh00, 8'sh20, 8'shfa, 8'shfb, 8'shec, 8'sh14
    /* (84, 0) */	    8'sh03, 8'shfc, 8'shf4, 8'sh07, 8'shfc, 8'sh19, 8'shf9, 8'shf7, 8'shfd, 8'sh03, 8'sh00, 8'sh1e, 8'shfb, 8'shfb, 8'shee, 8'sh13
    /* (85, 0) */	    8'sh03, 8'shfc, 8'shf5, 8'sh06, 8'shfc, 8'sh17, 8'shf9, 8'shf8, 8'shfd, 8'sh03, 8'sh00, 8'sh1b, 8'shfb, 8'shfc, 8'shef, 8'sh11
    /* (86, 0) */	    8'sh03, 8'shfc, 8'shf6, 8'sh06, 8'shfc, 8'sh15, 8'shfa, 8'shf9, 8'shfd, 8'sh02, 8'sh00, 8'sh19, 8'shfc, 8'shfc, 8'shf1, 8'sh0f
    /* (87, 0) */	    8'sh03, 8'shfd, 8'shf7, 8'sh05, 8'shfd, 8'sh13, 8'shfb, 8'shfa, 8'shfe, 8'sh02, 8'sh00, 8'sh16, 8'shfc, 8'shfc, 8'shf2, 8'sh0e
    /* (88, 0) */	    8'sh02, 8'shfd, 8'shf8, 8'sh05, 8'shfd, 8'sh11, 8'shfb, 8'shfa, 8'shfe, 8'sh02, 8'sh00, 8'sh14, 8'shfd, 8'shfd, 8'shf4, 8'sh0c
    /* (89, 0) */	    8'sh02, 8'shfd, 8'shf9, 8'sh04, 8'shfd, 8'sh0f, 8'shfc, 8'shfb, 8'shfe, 8'sh02, 8'sh00, 8'sh11, 8'shfd, 8'shfd, 8'shf5, 8'sh0b
    /* (90, 0) */	    8'sh02, 8'shfe, 8'shfa, 8'sh03, 8'shfe, 8'sh0d, 8'shfc, 8'shfc, 8'shfe, 8'sh01, 8'sh00, 8'sh0f, 8'shfd, 8'shfe, 8'shf7, 8'sh09
    /* (91, 0) */	    8'sh01, 8'shfe, 8'shfb, 8'sh03, 8'shfe, 8'sh0a, 8'shfd, 8'shfc, 8'shff, 8'sh01, 8'sh00, 8'sh0c, 8'shfe, 8'shfe, 8'shf8, 8'sh08
    /* (92, 0) */	    8'sh01, 8'shff, 8'shfc, 8'sh02, 8'shff, 8'sh08, 8'shfe, 8'shfd, 8'shff, 8'sh01, 8'sh00, 8'sh0a, 8'shfe, 8'shfe, 8'shfa, 8'sh06
    /* (93, 0) */	    8'sh01, 8'shff, 8'shfd, 8'sh02, 8'shff, 8'sh06, 8'shfe, 8'shfe, 8'shff, 8'sh01, 8'sh00, 8'sh07, 8'shff, 8'shff, 8'shfb, 8'sh05
    /* (94, 0) */	    8'sh01, 8'shff, 8'shfe, 8'sh01, 8'shff, 8'sh04, 8'shff, 8'shff, 8'shff, 8'sh00, 8'sh00, 8'sh05, 8'shff, 8'shff, 8'shfd, 8'sh03
    /* (95, 0) */	    8'sh00, 8'sh00, 8'shff, 8'sh01, 8'sh00, 8'sh02, 8'shff, 8'shff, 8'sh00, 8'sh00, 8'sh00, 8'sh02, 8'sh00, 8'sh00, 8'shfe, 8'sh02
    /* (96, 0) */	    8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00
    /* (97, 0) */	    8'sh00, 8'sh00, 8'sh01, 8'shff, 8'sh00, 8'shfe, 8'sh01, 8'sh01, 8'sh00, 8'sh00, 8'sh00, 8'shfe, 8'sh00, 8'sh00, 8'sh02, 8'shfe
    /* (98, 0) */	    8'shff, 8'sh01, 8'sh02, 8'shff, 8'sh01, 8'shfc, 8'sh01, 8'sh01, 8'sh01, 8'sh00, 8'sh00, 8'shfb, 8'sh01, 8'sh01, 8'sh03, 8'shfd
    /* (99, 0) */	    8'shff, 8'sh01, 8'sh03, 8'shfe, 8'sh01, 8'shfa, 8'sh02, 8'sh02, 8'sh01, 8'shff, 8'sh00, 8'shf9, 8'sh01, 8'sh01, 8'sh05, 8'shfb
    /* (100, 0) */	    8'shff, 8'sh01, 8'sh04, 8'shfe, 8'sh01, 8'shf8, 8'sh02, 8'sh03, 8'sh01, 8'shff, 8'sh00, 8'shf6, 8'sh02, 8'sh02, 8'sh06, 8'shfa
    /* (101, 0) */	    8'shff, 8'sh02, 8'sh05, 8'shfd, 8'sh02, 8'shf6, 8'sh03, 8'sh04, 8'sh01, 8'shff, 8'sh00, 8'shf4, 8'sh02, 8'sh02, 8'sh08, 8'shf8
    /* (102, 0) */	    8'shfe, 8'sh02, 8'sh06, 8'shfd, 8'sh02, 8'shf3, 8'sh04, 8'sh04, 8'sh02, 8'shff, 8'sh00, 8'shf1, 8'sh03, 8'sh02, 8'sh09, 8'shf7
    /* (103, 0) */	    8'shfe, 8'sh03, 8'sh07, 8'shfc, 8'sh03, 8'shf1, 8'sh04, 8'sh05, 8'sh02, 8'shfe, 8'sh00, 8'shef, 8'sh03, 8'sh03, 8'sh0b, 8'shf5
    /* (104, 0) */	    8'shfe, 8'sh03, 8'sh08, 8'shfb, 8'sh03, 8'shef, 8'sh05, 8'sh06, 8'sh02, 8'shfe, 8'sh00, 8'shec, 8'sh03, 8'sh03, 8'sh0c, 8'shf4
    /* (105, 0) */	    8'shfd, 8'sh03, 8'sh09, 8'shfb, 8'sh03, 8'shed, 8'sh05, 8'sh06, 8'sh02, 8'shfe, 8'sh00, 8'shea, 8'sh04, 8'sh04, 8'sh0e, 8'shf2
    /* (106, 0) */	    8'shfd, 8'sh04, 8'sh0a, 8'shfa, 8'sh04, 8'sheb, 8'sh06, 8'sh07, 8'sh03, 8'shfe, 8'sh00, 8'she7, 8'sh04, 8'sh04, 8'sh0f, 8'shf1
    /* (107, 0) */	    8'shfd, 8'sh04, 8'sh0b, 8'shfa, 8'sh04, 8'she9, 8'sh07, 8'sh08, 8'sh03, 8'shfd, 8'sh00, 8'she5, 8'sh05, 8'sh04, 8'sh11, 8'shef
    /* (108, 0) */	    8'shfd, 8'sh04, 8'sh0c, 8'shf9, 8'sh04, 8'she7, 8'sh07, 8'sh09, 8'sh03, 8'shfd, 8'sh00, 8'she2, 8'sh05, 8'sh05, 8'sh12, 8'shed
    /* (109, 0) */	    8'shfc, 8'sh05, 8'sh0d, 8'shf9, 8'sh05, 8'she5, 8'sh08, 8'sh09, 8'sh03, 8'shfd, 8'sh00, 8'she0, 8'sh06, 8'sh05, 8'sh14, 8'shec
    /* (110, 0) */	    8'shfc, 8'sh05, 8'sh0e, 8'shf8, 8'sh05, 8'she3, 8'sh09, 8'sh0a, 8'sh04, 8'shfd, 8'sh00, 8'shdd, 8'sh06, 8'sh06, 8'sh15, 8'shea
    /* (111, 0) */	    8'shfc, 8'sh06, 8'sh0f, 8'shf7, 8'sh05, 8'she1, 8'sh09, 8'sh0b, 8'sh04, 8'shfc, 8'sh00, 8'shdb, 8'sh07, 8'sh06, 8'sh17, 8'she9
    /* (112, 0) */	    8'shfb, 8'sh06, 8'sh10, 8'shf7, 8'sh06, 8'shde, 8'sh0a, 8'sh0b, 8'sh04, 8'shfc, 8'sh00, 8'shd8, 8'sh07, 8'sh06, 8'sh18, 8'she7
    /* (113, 0) */	    8'shfb, 8'sh06, 8'sh11, 8'shf6, 8'sh06, 8'shdc, 8'sh0a, 8'sh0c, 8'sh05, 8'shfc, 8'sh00, 8'shd6, 8'sh07, 8'sh07, 8'sh1a, 8'she6
    /* (114, 0) */	    8'shfb, 8'sh07, 8'sh12, 8'shf6, 8'sh06, 8'shda, 8'sh0b, 8'sh0d, 8'sh05, 8'shfc, 8'sh00, 8'shd3, 8'sh08, 8'sh07, 8'sh1b, 8'she4
    /* (115, 0) */	    8'shfb, 8'sh07, 8'sh13, 8'shf5, 8'sh07, 8'shd8, 8'sh0c, 8'sh0e, 8'sh05, 8'shfb, 8'sh00, 8'shd1, 8'sh08, 8'sh08, 8'sh1d, 8'she3
    /* (116, 0) */	    8'shfa, 8'sh07, 8'sh14, 8'shf5, 8'sh07, 8'shd6, 8'sh0c, 8'sh0e, 8'sh05, 8'shfb, 8'sh00, 8'shce, 8'sh09, 8'sh08, 8'sh1e, 8'she1
    /* (117, 0) */	    8'shfa, 8'sh08, 8'sh15, 8'shf4, 8'sh08, 8'shd4, 8'sh0d, 8'sh0f, 8'sh06, 8'shfb, 8'sh00, 8'shcc, 8'sh09, 8'sh08, 8'sh20, 8'shdf
    /* (118, 0) */	    8'shfa, 8'sh08, 8'sh16, 8'shf3, 8'sh08, 8'shd2, 8'sh0d, 8'sh10, 8'sh06, 8'shfb, 8'sh01, 8'shc9, 8'sh0a, 8'sh09, 8'sh21, 8'shde
    /* (119, 0) */	    8'shf9, 8'sh09, 8'sh17, 8'shf3, 8'sh08, 8'shd0, 8'sh0e, 8'sh10, 8'sh06, 8'shfa, 8'sh01, 8'shc7, 8'sh0a, 8'sh09, 8'sh23, 8'shdc
    /* (120, 0) */	    8'shf9, 8'sh09, 8'sh18, 8'shf2, 8'sh09, 8'shce, 8'sh0f, 8'sh11, 8'sh06, 8'shfa, 8'sh01, 8'shc4, 8'sh0a, 8'sh0a, 8'sh24, 8'shdb
    /* (121, 0) */	    8'shf9, 8'sh09, 8'sh19, 8'shf2, 8'sh09, 8'shcc, 8'sh0f, 8'sh12, 8'sh07, 8'shfa, 8'sh01, 8'shc2, 8'sh0b, 8'sh0a, 8'sh26, 8'shd9
    /* (122, 0) */	    8'shf9, 8'sh0a, 8'sh1a, 8'shf1, 8'sh09, 8'shca, 8'sh10, 8'sh13, 8'sh07, 8'shfa, 8'sh01, 8'shbf, 8'sh0b, 8'sh0a, 8'sh27, 8'shd8
    /* (123, 0) */	    8'shf8, 8'sh0a, 8'sh1b, 8'shf1, 8'sh0a, 8'shc7, 8'sh10, 8'sh13, 8'sh07, 8'shf9, 8'sh01, 8'shbd, 8'sh0c, 8'sh0b, 8'sh29, 8'shd6
    /* (124, 0) */	    8'shf8, 8'sh0a, 8'sh1c, 8'shf0, 8'sh0a, 8'shc5, 8'sh11, 8'sh14, 8'sh07, 8'shf9, 8'sh01, 8'shba, 8'sh0c, 8'sh0b, 8'sh2a, 8'shd5
    /* (125, 0) */	    8'shf8, 8'sh0b, 8'sh1d, 8'shef, 8'sh0a, 8'shc3, 8'sh12, 8'sh15, 8'sh08, 8'shf9, 8'sh01, 8'shb8, 8'sh0d, 8'sh0c, 8'sh2c, 8'shd3
    /* (126, 0) */	    8'shf7, 8'sh0b, 8'sh1e, 8'shef, 8'sh0b, 8'shc1, 8'sh12, 8'sh15, 8'sh08, 8'shf9, 8'sh01, 8'shb5, 8'sh0d, 8'sh0c, 8'sh2d, 8'shd2
    /* (127, 0) */	    8'shf7, 8'sh0c, 8'sh1f, 8'shee, 8'sh0b, 8'shbf, 8'sh13, 8'sh16, 8'sh08, 8'shf8, 8'sh01, 8'shb3, 8'sh0e, 8'sh0c, 8'sh2f, 8'shd0
    /* (128, 0) */	    8'shfa, 8'sh39, 8'shfb, 8'sh37, 8'shf6, 8'sh7f, 8'sh80, 8'sh38, 8'shed, 8'she4, 8'shf0, 8'shd6, 8'shc9, 8'sh12, 8'shda, 8'she2
    /* (129, 0) */	    8'shfa, 8'sh37, 8'shfb, 8'sh36, 8'shf6, 8'sh7b, 8'sh84, 8'sh36, 8'shee, 8'she5, 8'shf0, 8'shd7, 8'shcb, 8'sh11, 8'shdb, 8'she3
    /* (130, 0) */	    8'shfa, 8'sh35, 8'shfb, 8'sh34, 8'shf6, 8'sh78, 8'sh88, 8'sh34, 8'shee, 8'she6, 8'shf1, 8'shd9, 8'shcd, 8'sh11, 8'shdc, 8'she4
    /* (131, 0) */	    8'shfa, 8'sh33, 8'shfb, 8'sh32, 8'shf7, 8'sh74, 8'sh8c, 8'sh32, 8'shef, 8'she7, 8'shf1, 8'shda, 8'shce, 8'sh10, 8'shde, 8'she5
    /* (132, 0) */	    8'shfb, 8'sh32, 8'shfb, 8'sh30, 8'shf7, 8'sh70, 8'sh90, 8'sh31, 8'shef, 8'she8, 8'shf2, 8'shdb, 8'shd0, 8'sh10, 8'shdf, 8'she6
    /* (133, 0) */	    8'shfb, 8'sh30, 8'shfc, 8'sh2f, 8'shf7, 8'sh6c, 8'sh94, 8'sh2f, 8'shf0, 8'she9, 8'shf2, 8'shdd, 8'shd2, 8'sh0f, 8'she0, 8'she7
    /* (134, 0) */	    8'shfb, 8'sh2e, 8'shfc, 8'sh2d, 8'shf8, 8'sh68, 8'sh98, 8'sh2d, 8'shf1, 8'shea, 8'shf3, 8'shde, 8'shd3, 8'sh0e, 8'she1, 8'she8
    /* (135, 0) */	    8'shfb, 8'sh2c, 8'shfc, 8'sh2b, 8'shf8, 8'sh64, 8'sh9c, 8'sh2b, 8'shf1, 8'shea, 8'shf3, 8'shdf, 8'shd5, 8'sh0e, 8'she2, 8'she9
    /* (136, 0) */	    8'shfb, 8'sh2b, 8'shfc, 8'sh29, 8'shf8, 8'sh60, 8'sha0, 8'sh2a, 8'shf2, 8'sheb, 8'shf4, 8'she1, 8'shd7, 8'sh0d, 8'she4, 8'shea
    /* (137, 0) */	    8'shfc, 8'sh29, 8'shfc, 8'sh28, 8'shf9, 8'sh5c, 8'sha4, 8'sh28, 8'shf2, 8'shec, 8'shf4, 8'she2, 8'shd9, 8'sh0d, 8'she5, 8'sheb
    /* (138, 0) */	    8'shfc, 8'sh27, 8'shfc, 8'sh26, 8'shf9, 8'sh58, 8'sha8, 8'sh26, 8'shf3, 8'shed, 8'shf5, 8'she3, 8'shda, 8'sh0c, 8'she6, 8'shec
    /* (139, 0) */	    8'shfc, 8'sh25, 8'shfd, 8'sh24, 8'shf9, 8'sh54, 8'shac, 8'sh24, 8'shf4, 8'shee, 8'shf5, 8'she5, 8'shdc, 8'sh0c, 8'she7, 8'shed
    /* (140, 0) */	    8'shfc, 8'sh23, 8'shfd, 8'sh23, 8'shfa, 8'sh50, 8'shb0, 8'sh23, 8'shf4, 8'shef, 8'shf6, 8'she6, 8'shde, 8'sh0b, 8'she8, 8'shee
    /* (141, 0) */	    8'shfc, 8'sh22, 8'shfd, 8'sh21, 8'shfa, 8'sh4c, 8'shb4, 8'sh21, 8'shf5, 8'shf0, 8'shf6, 8'she7, 8'shdf, 8'sh0b, 8'shea, 8'shee
    /* (142, 0) */	    8'shfd, 8'sh20, 8'shfd, 8'sh1f, 8'shfa, 8'sh48, 8'shb8, 8'sh1f, 8'shf5, 8'shf0, 8'shf7, 8'she8, 8'she1, 8'sh0a, 8'sheb, 8'shef
    /* (143, 0) */	    8'shfd, 8'sh1e, 8'shfd, 8'sh1d, 8'shfb, 8'sh44, 8'shbc, 8'sh1e, 8'shf6, 8'shf1, 8'shf7, 8'shea, 8'she3, 8'sh09, 8'shec, 8'shf0
    /* (144, 0) */	    8'shfd, 8'sh1c, 8'shfd, 8'sh1c, 8'shfb, 8'sh40, 8'shc0, 8'sh1c, 8'shf7, 8'shf2, 8'shf8, 8'sheb, 8'she5, 8'sh09, 8'shed, 8'shf1
    /* (145, 0) */	    8'shfd, 8'sh1b, 8'shfe, 8'sh1a, 8'shfb, 8'sh3c, 8'shc4, 8'sh1a, 8'shf7, 8'shf3, 8'shf8, 8'shec, 8'she6, 8'sh08, 8'shee, 8'shf2
    /* (146, 0) */	    8'shfd, 8'sh19, 8'shfe, 8'sh18, 8'shfb, 8'sh38, 8'shc8, 8'sh18, 8'shf8, 8'shf4, 8'shf9, 8'shee, 8'she8, 8'sh08, 8'shef, 8'shf3
    /* (147, 0) */	    8'shfd, 8'sh17, 8'shfe, 8'sh16, 8'shfc, 8'sh34, 8'shcc, 8'sh17, 8'shf8, 8'shf5, 8'shf9, 8'shef, 8'shea, 8'sh07, 8'shf1, 8'shf4
    /* (148, 0) */	    8'shfe, 8'sh15, 8'shfe, 8'sh15, 8'shfc, 8'sh30, 8'shd0, 8'sh15, 8'shf9, 8'shf6, 8'shfa, 8'shf0, 8'sheb, 8'sh07, 8'shf2, 8'shf5
    /* (149, 0) */	    8'shfe, 8'sh13, 8'shfe, 8'sh13, 8'shfc, 8'sh2c, 8'shd4, 8'sh13, 8'shf9, 8'shf7, 8'shfa, 8'shf2, 8'shed, 8'sh06, 8'shf3, 8'shf6
    /* (150, 0) */	    8'shfe, 8'sh12, 8'shfe, 8'sh11, 8'shfd, 8'sh28, 8'shd8, 8'sh11, 8'shfa, 8'shf7, 8'shfb, 8'shf3, 8'shef, 8'sh06, 8'shf4, 8'shf7
    /* (151, 0) */	    8'shfe, 8'sh10, 8'shff, 8'sh10, 8'shfd, 8'sh24, 8'shdc, 8'sh10, 8'shfb, 8'shf8, 8'shfb, 8'shf4, 8'shf1, 8'sh05, 8'shf5, 8'shf8
    /* (152, 0) */	    8'shfe, 8'sh0e, 8'shff, 8'sh0e, 8'shfd, 8'sh20, 8'she0, 8'sh0e, 8'shfb, 8'shf9, 8'shfc, 8'shf6, 8'shf2, 8'sh04, 8'shf7, 8'shf9
    /* (153, 0) */	    8'shff, 8'sh0c, 8'shff, 8'sh0c, 8'shfe, 8'sh1c, 8'she4, 8'sh0c, 8'shfc, 8'shfa, 8'shfc, 8'shf7, 8'shf4, 8'sh04, 8'shf8, 8'shfa
    /* (154, 0) */	    8'shff, 8'sh0b, 8'shff, 8'sh0a, 8'shfe, 8'sh18, 8'she8, 8'sh0a, 8'shfc, 8'shfb, 8'shfd, 8'shf8, 8'shf6, 8'sh03, 8'shf9, 8'shfa
    /* (155, 0) */	    8'shff, 8'sh09, 8'shff, 8'sh09, 8'shfe, 8'sh14, 8'shec, 8'sh09, 8'shfd, 8'shfc, 8'shfd, 8'shf9, 8'shf7, 8'sh03, 8'shfa, 8'shfb
    /* (156, 0) */	    8'shff, 8'sh07, 8'shff, 8'sh07, 8'shff, 8'sh10, 8'shf0, 8'sh07, 8'shfe, 8'shfd, 8'shfe, 8'shfb, 8'shf9, 8'sh02, 8'shfb, 8'shfc
    /* (157, 0) */	    8'shff, 8'sh05, 8'sh00, 8'sh05, 8'shff, 8'sh0c, 8'shf4, 8'sh05, 8'shfe, 8'shfd, 8'shfe, 8'shfc, 8'shfb, 8'sh02, 8'shfc, 8'shfd
    /* (158, 0) */	    8'sh00, 8'sh04, 8'sh00, 8'sh03, 8'shff, 8'sh08, 8'shf8, 8'sh03, 8'shff, 8'shfe, 8'shff, 8'shfd, 8'shfd, 8'sh01, 8'shfe, 8'shfe
    /* (159, 0) */	    8'sh00, 8'sh02, 8'sh00, 8'sh02, 8'sh00, 8'sh04, 8'shfc, 8'sh02, 8'shff, 8'shff, 8'shff, 8'shff, 8'shfe, 8'sh01, 8'shff, 8'shff
    /* (160, 0) */	    8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00
    /* (161, 0) */	    8'sh00, 8'shfe, 8'sh00, 8'shfe, 8'sh00, 8'shfc, 8'sh04, 8'shfe, 8'sh01, 8'sh01, 8'sh01, 8'sh01, 8'sh02, 8'shff, 8'sh01, 8'sh01
    /* (162, 0) */	    8'sh00, 8'shfc, 8'sh00, 8'shfd, 8'sh01, 8'shf8, 8'sh08, 8'shfd, 8'sh01, 8'sh02, 8'sh01, 8'sh03, 8'sh03, 8'shff, 8'sh02, 8'sh02
    /* (163, 0) */	    8'sh01, 8'shfb, 8'sh00, 8'shfb, 8'sh01, 8'shf4, 8'sh0c, 8'shfb, 8'sh02, 8'sh03, 8'sh02, 8'sh04, 8'sh05, 8'shfe, 8'sh04, 8'sh03
    /* (164, 0) */	    8'sh01, 8'shf9, 8'sh01, 8'shf9, 8'sh01, 8'shf0, 8'sh10, 8'shf9, 8'sh02, 8'sh03, 8'sh02, 8'sh05, 8'sh07, 8'shfe, 8'sh05, 8'sh04
    /* (165, 0) */	    8'sh01, 8'shf7, 8'sh01, 8'shf7, 8'sh02, 8'shec, 8'sh14, 8'shf7, 8'sh03, 8'sh04, 8'sh03, 8'sh07, 8'sh09, 8'shfd, 8'sh06, 8'sh05
    /* (166, 0) */	    8'sh01, 8'shf5, 8'sh01, 8'shf6, 8'sh02, 8'she8, 8'sh18, 8'shf6, 8'sh04, 8'sh05, 8'sh03, 8'sh08, 8'sh0a, 8'shfd, 8'sh07, 8'sh06
    /* (167, 0) */	    8'sh01, 8'shf4, 8'sh01, 8'shf4, 8'sh02, 8'she4, 8'sh1c, 8'shf4, 8'sh04, 8'sh06, 8'sh04, 8'sh09, 8'sh0c, 8'shfc, 8'sh08, 8'sh06
    /* (168, 0) */	    8'sh02, 8'shf2, 8'sh01, 8'shf2, 8'sh03, 8'she0, 8'sh20, 8'shf2, 8'sh05, 8'sh07, 8'sh04, 8'sh0a, 8'sh0e, 8'shfc, 8'sh09, 8'sh07
    /* (169, 0) */	    8'sh02, 8'shf0, 8'sh01, 8'shf0, 8'sh03, 8'shdc, 8'sh24, 8'shf0, 8'sh05, 8'sh08, 8'sh05, 8'sh0c, 8'sh0f, 8'shfb, 8'sh0b, 8'sh08
    /* (170, 0) */	    8'sh02, 8'shee, 8'sh02, 8'shef, 8'sh03, 8'shd8, 8'sh28, 8'shef, 8'sh06, 8'sh09, 8'sh05, 8'sh0d, 8'sh11, 8'shfa, 8'sh0c, 8'sh09
    /* (171, 0) */	    8'sh02, 8'shed, 8'sh02, 8'shed, 8'sh04, 8'shd4, 8'sh2c, 8'shed, 8'sh07, 8'sh09, 8'sh06, 8'sh0e, 8'sh13, 8'shfa, 8'sh0d, 8'sh0a
    /* (172, 0) */	    8'sh02, 8'sheb, 8'sh02, 8'sheb, 8'sh04, 8'shd0, 8'sh30, 8'sheb, 8'sh07, 8'sh0a, 8'sh06, 8'sh10, 8'sh15, 8'shf9, 8'sh0e, 8'sh0b
    /* (173, 0) */	    8'sh03, 8'she9, 8'sh02, 8'shea, 8'sh04, 8'shcc, 8'sh34, 8'she9, 8'sh08, 8'sh0b, 8'sh07, 8'sh11, 8'sh16, 8'shf9, 8'sh0f, 8'sh0c
    /* (174, 0) */	    8'sh03, 8'she7, 8'sh02, 8'she8, 8'sh05, 8'shc8, 8'sh38, 8'she8, 8'sh08, 8'sh0c, 8'sh07, 8'sh12, 8'sh18, 8'shf8, 8'sh11, 8'sh0d
    /* (175, 0) */	    8'sh03, 8'she5, 8'sh02, 8'she6, 8'sh05, 8'shc4, 8'sh3c, 8'she6, 8'sh09, 8'sh0d, 8'sh08, 8'sh14, 8'sh1a, 8'shf8, 8'sh12, 8'sh0e
    /* (176, 0) */	    8'sh03, 8'she4, 8'sh03, 8'she4, 8'sh05, 8'shc0, 8'sh40, 8'she4, 8'sh09, 8'sh0e, 8'sh08, 8'sh15, 8'sh1b, 8'shf7, 8'sh13, 8'sh0f
    /* (177, 0) */	    8'sh03, 8'she2, 8'sh03, 8'she3, 8'sh05, 8'shbc, 8'sh44, 8'she2, 8'sh0a, 8'sh0f, 8'sh09, 8'sh16, 8'sh1d, 8'shf7, 8'sh14, 8'sh10
    /* (178, 0) */	    8'sh03, 8'she0, 8'sh03, 8'she1, 8'sh06, 8'shb8, 8'sh48, 8'she1, 8'sh0b, 8'sh10, 8'sh09, 8'sh18, 8'sh1f, 8'shf6, 8'sh15, 8'sh11
    /* (179, 0) */	    8'sh04, 8'shde, 8'sh03, 8'shdf, 8'sh06, 8'shb4, 8'sh4c, 8'shdf, 8'sh0b, 8'sh10, 8'sh0a, 8'sh19, 8'sh21, 8'shf5, 8'sh16, 8'sh12
    /* (180, 0) */	    8'sh04, 8'shdd, 8'sh03, 8'shdd, 8'sh06, 8'shb0, 8'sh50, 8'shdd, 8'sh0c, 8'sh11, 8'sh0a, 8'sh1a, 8'sh22, 8'shf5, 8'sh18, 8'sh12
    /* (181, 0) */	    8'sh04, 8'shdb, 8'sh03, 8'shdc, 8'sh07, 8'shac, 8'sh54, 8'shdc, 8'sh0c, 8'sh12, 8'sh0b, 8'sh1b, 8'sh24, 8'shf4, 8'sh19, 8'sh13
    /* (182, 0) */	    8'sh04, 8'shd9, 8'sh04, 8'shda, 8'sh07, 8'sha8, 8'sh58, 8'shda, 8'sh0d, 8'sh13, 8'sh0b, 8'sh1d, 8'sh26, 8'shf4, 8'sh1a, 8'sh14
    /* (183, 0) */	    8'sh04, 8'shd7, 8'sh04, 8'shd8, 8'sh07, 8'sha4, 8'sh5c, 8'shd8, 8'sh0e, 8'sh14, 8'sh0c, 8'sh1e, 8'sh27, 8'shf3, 8'sh1b, 8'sh15
    /* (184, 0) */	    8'sh05, 8'shd5, 8'sh04, 8'shd7, 8'sh08, 8'sha0, 8'sh60, 8'shd6, 8'sh0e, 8'sh15, 8'sh0c, 8'sh1f, 8'sh29, 8'shf3, 8'sh1c, 8'sh16
    /* (185, 0) */	    8'sh05, 8'shd4, 8'sh04, 8'shd5, 8'sh08, 8'sh9c, 8'sh64, 8'shd5, 8'sh0f, 8'sh16, 8'sh0d, 8'sh21, 8'sh2b, 8'shf2, 8'sh1e, 8'sh17
    /* (186, 0) */	    8'sh05, 8'shd2, 8'sh04, 8'shd3, 8'sh08, 8'sh98, 8'sh68, 8'shd3, 8'sh0f, 8'sh16, 8'sh0d, 8'sh22, 8'sh2d, 8'shf2, 8'sh1f, 8'sh18
    /* (187, 0) */	    8'sh05, 8'shd0, 8'sh04, 8'shd1, 8'sh09, 8'sh94, 8'sh6c, 8'shd1, 8'sh10, 8'sh17, 8'sh0e, 8'sh23, 8'sh2e, 8'shf1, 8'sh20, 8'sh19
    /* (188, 0) */	    8'sh05, 8'shce, 8'sh05, 8'shd0, 8'sh09, 8'sh90, 8'sh70, 8'shcf, 8'sh11, 8'sh18, 8'sh0e, 8'sh25, 8'sh30, 8'shf0, 8'sh21, 8'sh1a
    /* (189, 0) */	    8'sh06, 8'shcd, 8'sh05, 8'shce, 8'sh09, 8'sh8c, 8'sh74, 8'shce, 8'sh11, 8'sh19, 8'sh0f, 8'sh26, 8'sh32, 8'shf0, 8'sh22, 8'sh1b
    /* (190, 0) */	    8'sh06, 8'shcb, 8'sh05, 8'shcc, 8'sh0a, 8'sh88, 8'sh78, 8'shcc, 8'sh12, 8'sh1a, 8'sh0f, 8'sh27, 8'sh33, 8'shef, 8'sh24, 8'sh1c
    /* (191, 0) */	    8'sh06, 8'shc9, 8'sh05, 8'shca, 8'sh0a, 8'sh85, 8'sh7c, 8'shca, 8'sh12, 8'sh1b, 8'sh10, 8'sh29, 8'sh35, 8'shef, 8'sh25, 8'sh1d
    /* (192, 0) */	    8'sh2e, 8'shfb, 8'shf7, 8'she8, 8'shf4, 8'sh10, 8'sh0c, 8'sh18, 8'shf6, 8'sh23, 8'shfa, 8'sh15, 8'shff, 8'shff, 8'shd2, 8'shfc
    /* (193, 0) */	    8'sh2c, 8'shfb, 8'shf7, 8'she8, 8'shf5, 8'sh0f, 8'sh0c, 8'sh18, 8'shf6, 8'sh22, 8'shfb, 8'sh14, 8'shff, 8'shff, 8'shd3, 8'shfc
    /* (194, 0) */	    8'sh2b, 8'shfb, 8'shf8, 8'she9, 8'shf5, 8'sh0f, 8'sh0b, 8'sh17, 8'shf6, 8'sh21, 8'shfb, 8'sh14, 8'shff, 8'shff, 8'shd5, 8'shfd
    /* (195, 0) */	    8'sh2a, 8'shfb, 8'shf8, 8'shea, 8'shf5, 8'sh0e, 8'sh0b, 8'sh16, 8'shf7, 8'sh20, 8'shfb, 8'sh13, 8'sh00, 8'shff, 8'shd6, 8'shfd
    /* (196, 0) */	    8'sh28, 8'shfb, 8'shf8, 8'sheb, 8'shf6, 8'sh0e, 8'sh0b, 8'sh15, 8'shf7, 8'sh1f, 8'shfb, 8'sh12, 8'sh00, 8'shff, 8'shd8, 8'shfd
    /* (197, 0) */	    8'sh27, 8'shfc, 8'shf8, 8'sheb, 8'shf6, 8'sh0d, 8'sh0a, 8'sh14, 8'shf7, 8'sh1e, 8'shfb, 8'sh12, 8'sh00, 8'shff, 8'shd9, 8'shfd
    /* (198, 0) */	    8'sh25, 8'shfc, 8'shf9, 8'shec, 8'shf6, 8'sh0d, 8'sh0a, 8'sh14, 8'shf8, 8'sh1d, 8'shfb, 8'sh11, 8'sh00, 8'shff, 8'shda, 8'shfd
    /* (199, 0) */	    8'sh24, 8'shfc, 8'shf9, 8'shed, 8'shf7, 8'sh0c, 8'sh09, 8'sh13, 8'shf8, 8'sh1c, 8'shfc, 8'sh10, 8'sh00, 8'shff, 8'shdc, 8'shfd
    /* (200, 0) */	    8'sh22, 8'shfc, 8'shf9, 8'shee, 8'shf7, 8'sh0c, 8'sh09, 8'sh12, 8'shf8, 8'sh1b, 8'shfc, 8'sh10, 8'sh00, 8'shff, 8'shdd, 8'shfd
    /* (201, 0) */	    8'sh21, 8'shfc, 8'shfa, 8'shef, 8'shf8, 8'sh0b, 8'sh09, 8'sh11, 8'shf9, 8'sh19, 8'shfc, 8'sh0f, 8'sh00, 8'shff, 8'shdf, 8'shfd
    /* (202, 0) */	    8'sh1f, 8'shfc, 8'shfa, 8'shef, 8'shf8, 8'sh0b, 8'sh08, 8'sh11, 8'shf9, 8'sh18, 8'shfc, 8'sh0e, 8'sh00, 8'shff, 8'she0, 8'shfd
    /* (203, 0) */	    8'sh1e, 8'shfd, 8'shfa, 8'shf0, 8'shf8, 8'sh0a, 8'sh08, 8'sh10, 8'shf9, 8'sh17, 8'shfc, 8'sh0e, 8'sh00, 8'shff, 8'she2, 8'shfe
    /* (204, 0) */	    8'sh1d, 8'shfd, 8'shfa, 8'shf1, 8'shf9, 8'sh0a, 8'sh08, 8'sh0f, 8'shfa, 8'sh16, 8'shfd, 8'sh0d, 8'sh00, 8'shff, 8'she3, 8'shfe
    /* (205, 0) */	    8'sh1b, 8'shfd, 8'shfb, 8'shf2, 8'shf9, 8'sh09, 8'sh07, 8'sh0e, 8'shfa, 8'sh15, 8'shfd, 8'sh0c, 8'sh00, 8'shff, 8'she5, 8'shfe
    /* (206, 0) */	    8'sh1a, 8'shfd, 8'shfb, 8'shf2, 8'shf9, 8'sh09, 8'sh07, 8'sh0e, 8'shfa, 8'sh14, 8'shfd, 8'sh0c, 8'sh00, 8'shff, 8'she6, 8'shfe
    /* (207, 0) */	    8'sh18, 8'shfd, 8'shfb, 8'shf3, 8'shfa, 8'sh08, 8'sh06, 8'sh0d, 8'shfb, 8'sh13, 8'shfd, 8'sh0b, 8'sh00, 8'shff, 8'she7, 8'shfe
    /* (208, 0) */	    8'sh17, 8'shfd, 8'shfb, 8'shf4, 8'shfa, 8'sh08, 8'sh06, 8'sh0c, 8'shfb, 8'sh12, 8'shfd, 8'sh0a, 8'sh00, 8'shff, 8'she9, 8'shfe
    /* (209, 0) */	    8'sh15, 8'shfe, 8'shfc, 8'shf5, 8'shfa, 8'sh07, 8'sh06, 8'sh0b, 8'shfb, 8'sh11, 8'shfd, 8'sh0a, 8'sh00, 8'shff, 8'shea, 8'shfe
    /* (210, 0) */	    8'sh14, 8'shfe, 8'shfc, 8'shf5, 8'shfb, 8'sh07, 8'sh05, 8'sh0b, 8'shfc, 8'sh0f, 8'shfe, 8'sh09, 8'sh00, 8'shff, 8'shec, 8'shfe
    /* (211, 0) */	    8'sh13, 8'shfe, 8'shfc, 8'shf6, 8'shfb, 8'sh06, 8'sh05, 8'sh0a, 8'shfc, 8'sh0e, 8'shfe, 8'sh08, 8'sh00, 8'sh00, 8'shed, 8'shfe
    /* (212, 0) */	    8'sh11, 8'shfe, 8'shfd, 8'shf7, 8'shfc, 8'sh06, 8'sh05, 8'sh09, 8'shfc, 8'sh0d, 8'shfe, 8'sh08, 8'sh00, 8'sh00, 8'shef, 8'shff
    /* (213, 0) */	    8'sh10, 8'shfe, 8'shfd, 8'shf8, 8'shfc, 8'sh05, 8'sh04, 8'sh08, 8'shfc, 8'sh0c, 8'shfe, 8'sh07, 8'sh00, 8'sh00, 8'shf0, 8'shff
    /* (214, 0) */	    8'sh0e, 8'shfe, 8'shfd, 8'shf8, 8'shfc, 8'sh05, 8'sh04, 8'sh08, 8'shfd, 8'sh0b, 8'shfe, 8'sh07, 8'sh00, 8'sh00, 8'shf2, 8'shff
    /* (215, 0) */	    8'sh0d, 8'shff, 8'shfd, 8'shf9, 8'shfd, 8'sh04, 8'sh03, 8'sh07, 8'shfd, 8'sh0a, 8'shfe, 8'sh06, 8'sh00, 8'sh00, 8'shf3, 8'shff
    /* (216, 0) */	    8'sh0b, 8'shff, 8'shfe, 8'shfa, 8'shfd, 8'sh04, 8'sh03, 8'sh06, 8'shfd, 8'sh09, 8'shff, 8'sh05, 8'sh00, 8'sh00, 8'shf4, 8'shff
    /* (217, 0) */	    8'sh0a, 8'shff, 8'shfe, 8'shfb, 8'shfd, 8'sh03, 8'sh03, 8'sh05, 8'shfe, 8'sh08, 8'shff, 8'sh05, 8'sh00, 8'sh00, 8'shf6, 8'shff
    /* (218, 0) */	    8'sh09, 8'shff, 8'shfe, 8'shfb, 8'shfe, 8'sh03, 8'sh02, 8'sh05, 8'shfe, 8'sh07, 8'shff, 8'sh04, 8'sh00, 8'sh00, 8'shf7, 8'shff
    /* (219, 0) */	    8'sh07, 8'shff, 8'shff, 8'shfc, 8'shfe, 8'sh02, 8'sh02, 8'sh04, 8'shfe, 8'sh06, 8'shff, 8'sh03, 8'sh00, 8'sh00, 8'shf9, 8'shff
    /* (220, 0) */	    8'sh06, 8'shff, 8'shff, 8'shfd, 8'shff, 8'sh02, 8'sh02, 8'sh03, 8'shff, 8'sh04, 8'shff, 8'sh03, 8'sh00, 8'sh00, 8'shfa, 8'sh00
    /* (221, 0) */	    8'sh04, 8'sh00, 8'shff, 8'shfe, 8'shff, 8'sh01, 8'sh01, 8'sh02, 8'shff, 8'sh03, 8'shff, 8'sh02, 8'sh00, 8'sh00, 8'shfc, 8'sh00
    /* (222, 0) */	    8'sh03, 8'sh00, 8'shff, 8'shfe, 8'shff, 8'sh01, 8'sh01, 8'sh02, 8'shff, 8'sh02, 8'sh00, 8'sh01, 8'sh00, 8'sh00, 8'shfd, 8'sh00
    /* (223, 0) */	    8'sh01, 8'sh00, 8'sh00, 8'shff, 8'sh00, 8'sh00, 8'sh00, 8'sh01, 8'sh00, 8'sh01, 8'sh00, 8'sh01, 8'sh00, 8'sh00, 8'shff, 8'sh00
    /* (224, 0) */	    8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00
    /* (225, 0) */	    8'shff, 8'sh00, 8'sh00, 8'sh01, 8'sh00, 8'sh00, 8'sh00, 8'shff, 8'sh00, 8'shff, 8'sh00, 8'shff, 8'sh00, 8'sh00, 8'sh01, 8'sh00
    /* (226, 0) */	    8'shfd, 8'sh00, 8'sh01, 8'sh02, 8'sh01, 8'shff, 8'shff, 8'shfe, 8'sh01, 8'shfe, 8'sh00, 8'shff, 8'sh00, 8'sh00, 8'sh03, 8'sh00
    /* (227, 0) */	    8'shfc, 8'sh00, 8'sh01, 8'sh02, 8'sh01, 8'shff, 8'shff, 8'shfe, 8'sh01, 8'shfd, 8'sh01, 8'shfe, 8'sh00, 8'sh00, 8'sh04, 8'sh00
    /* (228, 0) */	    8'shfa, 8'sh01, 8'sh01, 8'sh03, 8'sh01, 8'shfe, 8'shfe, 8'shfd, 8'sh01, 8'shfc, 8'sh01, 8'shfd, 8'sh00, 8'sh00, 8'sh06, 8'sh00
    /* (229, 0) */	    8'shf9, 8'sh01, 8'sh01, 8'sh04, 8'sh02, 8'shfe, 8'shfe, 8'shfc, 8'sh02, 8'shfa, 8'sh01, 8'shfd, 8'sh00, 8'sh00, 8'sh07, 8'sh01
    /* (230, 0) */	    8'shf7, 8'sh01, 8'sh02, 8'sh05, 8'sh02, 8'shfd, 8'shfe, 8'shfb, 8'sh02, 8'shf9, 8'sh01, 8'shfc, 8'sh00, 8'sh00, 8'sh09, 8'sh01
    /* (231, 0) */	    8'shf6, 8'sh01, 8'sh02, 8'sh05, 8'sh03, 8'shfd, 8'shfd, 8'shfb, 8'sh02, 8'shf8, 8'sh01, 8'shfb, 8'sh00, 8'sh00, 8'sh0a, 8'sh01
    /* (232, 0) */	    8'shf5, 8'sh01, 8'sh02, 8'sh06, 8'sh03, 8'shfc, 8'shfd, 8'shfa, 8'sh03, 8'shf7, 8'sh01, 8'shfb, 8'sh00, 8'sh00, 8'sh0c, 8'sh01
    /* (233, 0) */	    8'shf3, 8'sh01, 8'sh03, 8'sh07, 8'sh03, 8'shfc, 8'shfd, 8'shf9, 8'sh03, 8'shf6, 8'sh02, 8'shfa, 8'sh00, 8'sh00, 8'sh0d, 8'sh01
    /* (234, 0) */	    8'shf2, 8'sh02, 8'sh03, 8'sh08, 8'sh04, 8'shfb, 8'shfc, 8'shf8, 8'sh03, 8'shf5, 8'sh02, 8'shf9, 8'sh00, 8'sh00, 8'sh0e, 8'sh01
    /* (235, 0) */	    8'shf0, 8'sh02, 8'sh03, 8'sh08, 8'sh04, 8'shfb, 8'shfc, 8'shf8, 8'sh04, 8'shf4, 8'sh02, 8'shf9, 8'sh00, 8'sh00, 8'sh10, 8'sh01
    /* (236, 0) */	    8'shef, 8'sh02, 8'sh03, 8'sh09, 8'sh04, 8'shfa, 8'shfb, 8'shf7, 8'sh04, 8'shf3, 8'sh02, 8'shf8, 8'sh00, 8'sh00, 8'sh11, 8'sh01
    /* (237, 0) */	    8'shed, 8'sh02, 8'sh04, 8'sh0a, 8'sh05, 8'shfa, 8'shfb, 8'shf6, 8'sh04, 8'shf2, 8'sh02, 8'shf8, 8'sh00, 8'sh00, 8'sh13, 8'sh02
    /* (238, 0) */	    8'shec, 8'sh02, 8'sh04, 8'sh0b, 8'sh05, 8'shf9, 8'shfb, 8'shf5, 8'sh04, 8'shf1, 8'sh02, 8'shf7, 8'sh00, 8'sh01, 8'sh14, 8'sh02
    /* (239, 0) */	    8'sheb, 8'sh02, 8'sh04, 8'sh0b, 8'sh06, 8'shf9, 8'shfa, 8'shf5, 8'sh05, 8'shef, 8'sh03, 8'shf6, 8'sh00, 8'sh01, 8'sh16, 8'sh02
    /* (240, 0) */	    8'she9, 8'sh03, 8'sh05, 8'sh0c, 8'sh06, 8'shf8, 8'shfa, 8'shf4, 8'sh05, 8'shee, 8'sh03, 8'shf6, 8'sh00, 8'sh01, 8'sh17, 8'sh02
    /* (241, 0) */	    8'she8, 8'sh03, 8'sh05, 8'sh0d, 8'sh06, 8'shf8, 8'shfa, 8'shf3, 8'sh05, 8'shed, 8'sh03, 8'shf5, 8'sh00, 8'sh01, 8'sh19, 8'sh02
    /* (242, 0) */	    8'she6, 8'sh03, 8'sh05, 8'sh0e, 8'sh07, 8'shf7, 8'shf9, 8'shf2, 8'sh06, 8'shec, 8'sh03, 8'shf4, 8'sh00, 8'sh01, 8'sh1a, 8'sh02
    /* (243, 0) */	    8'she5, 8'sh03, 8'sh05, 8'sh0e, 8'sh07, 8'shf7, 8'shf9, 8'shf2, 8'sh06, 8'sheb, 8'sh03, 8'shf4, 8'sh00, 8'sh01, 8'sh1b, 8'sh02
    /* (244, 0) */	    8'she3, 8'sh03, 8'sh06, 8'sh0f, 8'sh07, 8'shf6, 8'shf8, 8'shf1, 8'sh06, 8'shea, 8'sh03, 8'shf3, 8'sh00, 8'sh01, 8'sh1d, 8'sh02
    /* (245, 0) */	    8'she2, 8'sh03, 8'sh06, 8'sh10, 8'sh08, 8'shf6, 8'shf8, 8'shf0, 8'sh07, 8'she9, 8'sh04, 8'shf2, 8'sh00, 8'sh01, 8'sh1e, 8'sh02
    /* (246, 0) */	    8'she1, 8'sh04, 8'sh06, 8'sh11, 8'sh08, 8'shf5, 8'shf8, 8'shef, 8'sh07, 8'she8, 8'sh04, 8'shf2, 8'sh00, 8'sh01, 8'sh20, 8'sh03
    /* (247, 0) */	    8'shdf, 8'sh04, 8'sh06, 8'sh11, 8'sh08, 8'shf5, 8'shf7, 8'shef, 8'sh07, 8'she7, 8'sh04, 8'shf1, 8'sh00, 8'sh01, 8'sh21, 8'sh03
    /* (248, 0) */	    8'shde, 8'sh04, 8'sh07, 8'sh12, 8'sh09, 8'shf4, 8'shf7, 8'shee, 8'sh08, 8'she5, 8'sh04, 8'shf0, 8'sh00, 8'sh01, 8'sh23, 8'sh03
    /* (249, 0) */	    8'shdc, 8'sh04, 8'sh07, 8'sh13, 8'sh09, 8'shf4, 8'shf7, 8'shed, 8'sh08, 8'she4, 8'sh04, 8'shf0, 8'sh00, 8'sh01, 8'sh24, 8'sh03
    /* (250, 0) */	    8'shdb, 8'sh04, 8'sh07, 8'sh14, 8'sh0a, 8'shf3, 8'shf6, 8'shec, 8'sh08, 8'she3, 8'sh05, 8'shef, 8'sh00, 8'sh01, 8'sh26, 8'sh03
    /* (251, 0) */	    8'shd9, 8'sh04, 8'sh08, 8'sh15, 8'sh0a, 8'shf3, 8'shf6, 8'shec, 8'sh09, 8'she2, 8'sh05, 8'shee, 8'sh00, 8'sh01, 8'sh27, 8'sh03
    /* (252, 0) */	    8'shd8, 8'sh05, 8'sh08, 8'sh15, 8'sh0a, 8'shf2, 8'shf5, 8'sheb, 8'sh09, 8'she1, 8'sh05, 8'shee, 8'sh00, 8'sh01, 8'sh28, 8'sh03
    /* (253, 0) */	    8'shd6, 8'sh05, 8'sh08, 8'sh16, 8'sh0b, 8'shf2, 8'shf5, 8'shea, 8'sh09, 8'she0, 8'sh05, 8'shed, 8'sh00, 8'sh01, 8'sh2a, 8'sh03
    /* (254, 0) */	    8'shd5, 8'sh05, 8'sh08, 8'sh17, 8'sh0b, 8'shf1, 8'shf5, 8'she9, 8'sh0a, 8'shdf, 8'sh05, 8'shec, 8'sh01, 8'sh01, 8'sh2b, 8'sh03
    /* (255, 0) */	    8'shd4, 8'sh05, 8'sh09, 8'sh18, 8'sh0b, 8'shf1, 8'shf4, 8'she8, 8'sh0a, 8'shde, 8'sh05, 8'shec, 8'sh01, 8'sh01, 8'sh2d, 8'sh04
    /* (256, 0) */	    8'shcf, 8'shcf, 8'sh7f, 8'sh7f, 8'shb7, 8'sha3, 8'shde, 8'shfe, 8'shb2, 8'shd1, 8'sh01, 8'sh9f, 8'sh7f, 8'sh33, 8'sh07, 8'shcf
    /* (257, 0) */	    8'shd1, 8'shd1, 8'sh7b, 8'sh7f, 8'shb9, 8'sha6, 8'shdf, 8'shfe, 8'shb4, 8'shd3, 8'sh01, 8'sha2, 8'sh7c, 8'sh31, 8'sh06, 8'shd0
    /* (258, 0) */	    8'shd2, 8'shd2, 8'sh77, 8'sh7f, 8'shbb, 8'sha9, 8'she0, 8'shff, 8'shb7, 8'shd4, 8'sh01, 8'sha5, 8'sh78, 8'sh30, 8'sh06, 8'shd2
    /* (259, 0) */	    8'shd4, 8'shd4, 8'sh74, 8'sh7c, 8'shbe, 8'shac, 8'she1, 8'shff, 8'shb9, 8'shd6, 8'sh01, 8'sha8, 8'sh74, 8'sh2e, 8'sh06, 8'shd3
    /* (260, 0) */	    8'shd5, 8'shd5, 8'sh70, 8'sh78, 8'shc0, 8'shae, 8'she2, 8'shff, 8'shbc, 8'shd7, 8'sh01, 8'shab, 8'sh70, 8'sh2d, 8'sh06, 8'shd5
    /* (261, 0) */	    8'shd7, 8'shd7, 8'sh6c, 8'sh74, 8'shc2, 8'shb1, 8'she3, 8'shff, 8'shbe, 8'shd9, 8'sh01, 8'shae, 8'sh6c, 8'sh2b, 8'sh06, 8'shd6
    /* (262, 0) */	    8'shd8, 8'shd8, 8'sh68, 8'sh6f, 8'shc5, 8'shb4, 8'she4, 8'shff, 8'shc1, 8'shda, 8'sh01, 8'shb1, 8'sh68, 8'sh29, 8'sh05, 8'shd8
    /* (263, 0) */	    8'shda, 8'shda, 8'sh64, 8'sh6b, 8'shc7, 8'shb7, 8'she5, 8'shff, 8'shc3, 8'shdc, 8'sh01, 8'shb4, 8'sh64, 8'sh28, 8'sh05, 8'shd9
    /* (264, 0) */	    8'shdb, 8'shdb, 8'sh60, 8'sh67, 8'shc9, 8'shba, 8'she6, 8'shff, 8'shc6, 8'shdd, 8'sh01, 8'shb7, 8'sh60, 8'sh26, 8'sh05, 8'shdb
    /* (265, 0) */	    8'shdd, 8'shdd, 8'sh5c, 8'sh63, 8'shcb, 8'shbd, 8'she8, 8'shff, 8'shc8, 8'shde, 8'sh01, 8'shba, 8'sh5c, 8'sh25, 8'sh05, 8'shdd
    /* (266, 0) */	    8'shde, 8'shde, 8'sh58, 8'sh5e, 8'shce, 8'shc0, 8'she9, 8'shff, 8'shca, 8'she0, 8'sh01, 8'shbd, 8'sh58, 8'sh23, 8'sh05, 8'shde
    /* (267, 0) */	    8'she0, 8'she0, 8'sh54, 8'sh5a, 8'shd0, 8'shc3, 8'shea, 8'shff, 8'shcd, 8'she1, 8'sh01, 8'shc1, 8'sh54, 8'sh21, 8'sh04, 8'she0
    /* (268, 0) */	    8'she1, 8'she1, 8'sh50, 8'sh56, 8'shd2, 8'shc6, 8'sheb, 8'shff, 8'shcf, 8'she3, 8'sh01, 8'shc4, 8'sh50, 8'sh20, 8'sh04, 8'she1
    /* (269, 0) */	    8'she3, 8'she3, 8'sh4c, 8'sh51, 8'shd5, 8'shc9, 8'shec, 8'shff, 8'shd2, 8'she4, 8'sh01, 8'shc7, 8'sh4c, 8'sh1e, 8'sh04, 8'she3
    /* (270, 0) */	    8'she5, 8'she5, 8'sh48, 8'sh4d, 8'shd7, 8'shcc, 8'shed, 8'shff, 8'shd4, 8'she6, 8'sh01, 8'shca, 8'sh48, 8'sh1d, 8'sh04, 8'she4
    /* (271, 0) */	    8'she6, 8'she6, 8'sh44, 8'sh49, 8'shd9, 8'shce, 8'shee, 8'shff, 8'shd7, 8'she7, 8'sh01, 8'shcd, 8'sh44, 8'sh1b, 8'sh04, 8'she6
    /* (272, 0) */	    8'she8, 8'she8, 8'sh40, 8'sh45, 8'shdb, 8'shd1, 8'shef, 8'shff, 8'shd9, 8'she9, 8'sh01, 8'shd0, 8'sh40, 8'sh19, 8'sh03, 8'she7
    /* (273, 0) */	    8'she9, 8'she9, 8'sh3c, 8'sh40, 8'shde, 8'shd4, 8'shf0, 8'shff, 8'shdb, 8'shea, 8'sh01, 8'shd3, 8'sh3c, 8'sh18, 8'sh03, 8'she9
    /* (274, 0) */	    8'sheb, 8'sheb, 8'sh38, 8'sh3c, 8'she0, 8'shd7, 8'shf1, 8'shff, 8'shde, 8'shec, 8'sh01, 8'shd6, 8'sh38, 8'sh16, 8'sh03, 8'shea
    /* (275, 0) */	    8'shec, 8'shec, 8'sh34, 8'sh38, 8'she2, 8'shda, 8'shf2, 8'shff, 8'she0, 8'shed, 8'sh01, 8'shd9, 8'sh34, 8'sh15, 8'sh03, 8'shec
    /* (276, 0) */	    8'shee, 8'shee, 8'sh30, 8'sh33, 8'she5, 8'shdd, 8'shf3, 8'shff, 8'she3, 8'shee, 8'sh01, 8'shdc, 8'sh30, 8'sh13, 8'sh02, 8'shee
    /* (277, 0) */	    8'shef, 8'shef, 8'sh2c, 8'sh2f, 8'she7, 8'she0, 8'shf4, 8'shff, 8'she5, 8'shf0, 8'sh01, 8'shdf, 8'sh2c, 8'sh12, 8'sh02, 8'shef
    /* (278, 0) */	    8'shf1, 8'shf1, 8'sh28, 8'sh2b, 8'she9, 8'she3, 8'shf5, 8'sh00, 8'she8, 8'shf1, 8'sh00, 8'she2, 8'sh28, 8'sh10, 8'sh02, 8'shf1
    /* (279, 0) */	    8'shf2, 8'shf2, 8'sh24, 8'sh27, 8'sheb, 8'she6, 8'shf6, 8'sh00, 8'shea, 8'shf3, 8'sh00, 8'she5, 8'sh24, 8'sh0e, 8'sh02, 8'shf2
    /* (280, 0) */	    8'shf4, 8'shf4, 8'sh20, 8'sh22, 8'shee, 8'she9, 8'shf7, 8'sh00, 8'shed, 8'shf4, 8'sh00, 8'she8, 8'sh20, 8'sh0d, 8'sh02, 8'shf4
    /* (281, 0) */	    8'shf5, 8'shf5, 8'sh1c, 8'sh1e, 8'shf0, 8'shec, 8'shf9, 8'sh00, 8'shef, 8'shf6, 8'sh00, 8'sheb, 8'sh1c, 8'sh0b, 8'sh01, 8'shf5
    /* (282, 0) */	    8'shf7, 8'shf7, 8'sh18, 8'sh1a, 8'shf2, 8'shef, 8'shfa, 8'sh00, 8'shf1, 8'shf7, 8'sh00, 8'shee, 8'sh18, 8'sh0a, 8'sh01, 8'shf7
    /* (283, 0) */	    8'shf8, 8'shf8, 8'sh14, 8'sh15, 8'shf5, 8'shf1, 8'shfb, 8'sh00, 8'shf4, 8'shf9, 8'sh00, 8'shf1, 8'sh14, 8'sh08, 8'sh01, 8'shf8
    /* (284, 0) */	    8'shfa, 8'shfa, 8'sh10, 8'sh11, 8'shf7, 8'shf4, 8'shfc, 8'sh00, 8'shf6, 8'shfa, 8'sh00, 8'shf4, 8'sh10, 8'sh06, 8'sh01, 8'shfa
    /* (285, 0) */	    8'shfb, 8'shfb, 8'sh0c, 8'sh0d, 8'shf9, 8'shf7, 8'shfd, 8'sh00, 8'shf9, 8'shfc, 8'sh00, 8'shf7, 8'sh0c, 8'sh05, 8'sh01, 8'shfb
    /* (286, 0) */	    8'shfd, 8'shfd, 8'sh08, 8'sh09, 8'shfb, 8'shfa, 8'shfe, 8'sh00, 8'shfb, 8'shfd, 8'sh00, 8'shfa, 8'sh08, 8'sh03, 8'sh00, 8'shfd
    /* (287, 0) */	    8'shfe, 8'shfe, 8'sh04, 8'sh04, 8'shfe, 8'shfd, 8'shff, 8'sh00, 8'shfe, 8'shff, 8'sh00, 8'shfd, 8'sh04, 8'sh02, 8'sh00, 8'shfe
    /* (288, 0) */	    8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00
    /* (289, 0) */	    8'sh02, 8'sh02, 8'shfc, 8'shfc, 8'sh02, 8'sh03, 8'sh01, 8'sh00, 8'sh02, 8'sh01, 8'sh00, 8'sh03, 8'shfc, 8'shfe, 8'sh00, 8'sh02
    /* (290, 0) */	    8'sh03, 8'sh03, 8'shf8, 8'shf7, 8'sh05, 8'sh06, 8'sh02, 8'sh00, 8'sh05, 8'sh03, 8'sh00, 8'sh06, 8'shf8, 8'shfd, 8'sh00, 8'sh03
    /* (291, 0) */	    8'sh05, 8'sh05, 8'shf4, 8'shf3, 8'sh07, 8'sh09, 8'sh03, 8'sh00, 8'sh07, 8'sh04, 8'sh00, 8'sh09, 8'shf4, 8'shfb, 8'shff, 8'sh05
    /* (292, 0) */	    8'sh06, 8'sh06, 8'shf0, 8'shef, 8'sh09, 8'sh0c, 8'sh04, 8'sh00, 8'sh0a, 8'sh06, 8'sh00, 8'sh0c, 8'shf0, 8'shfa, 8'shff, 8'sh06
    /* (293, 0) */	    8'sh08, 8'sh08, 8'shec, 8'sheb, 8'sh0b, 8'sh0f, 8'sh05, 8'sh00, 8'sh0c, 8'sh07, 8'sh00, 8'sh0f, 8'shec, 8'shf8, 8'shff, 8'sh08
    /* (294, 0) */	    8'sh09, 8'sh09, 8'she8, 8'she6, 8'sh0e, 8'sh11, 8'sh06, 8'sh00, 8'sh0f, 8'sh09, 8'sh00, 8'sh12, 8'she8, 8'shf6, 8'shff, 8'sh09
    /* (295, 0) */	    8'sh0b, 8'sh0b, 8'she4, 8'she2, 8'sh10, 8'sh14, 8'sh07, 8'sh00, 8'sh11, 8'sh0a, 8'sh00, 8'sh15, 8'she4, 8'shf5, 8'shff, 8'sh0b
    /* (296, 0) */	    8'sh0c, 8'sh0c, 8'she0, 8'shde, 8'sh12, 8'sh17, 8'sh09, 8'sh00, 8'sh13, 8'sh0c, 8'sh00, 8'sh18, 8'she0, 8'shf3, 8'shfe, 8'sh0c
    /* (297, 0) */	    8'sh0e, 8'sh0e, 8'shdc, 8'shd9, 8'sh15, 8'sh1a, 8'sh0a, 8'sh00, 8'sh16, 8'sh0d, 8'sh00, 8'sh1b, 8'shdc, 8'shf2, 8'shfe, 8'sh0e
    /* (298, 0) */	    8'sh0f, 8'sh0f, 8'shd8, 8'shd5, 8'sh17, 8'sh1d, 8'sh0b, 8'sh00, 8'sh18, 8'sh0f, 8'sh00, 8'sh1e, 8'shd8, 8'shf0, 8'shfe, 8'sh0f
    /* (299, 0) */	    8'sh11, 8'sh11, 8'shd4, 8'shd1, 8'sh19, 8'sh20, 8'sh0c, 8'sh01, 8'sh1b, 8'sh10, 8'shff, 8'sh21, 8'shd4, 8'shee, 8'shfe, 8'sh11
    /* (300, 0) */	    8'sh12, 8'sh12, 8'shd0, 8'shcd, 8'sh1b, 8'sh23, 8'sh0d, 8'sh01, 8'sh1d, 8'sh12, 8'shff, 8'sh24, 8'shd0, 8'shed, 8'shfe, 8'sh12
    /* (301, 0) */	    8'sh14, 8'sh14, 8'shcc, 8'shc8, 8'sh1e, 8'sh26, 8'sh0e, 8'sh01, 8'sh20, 8'sh13, 8'shff, 8'sh27, 8'shcc, 8'sheb, 8'shfd, 8'sh14
    /* (302, 0) */	    8'sh15, 8'sh15, 8'shc8, 8'shc4, 8'sh20, 8'sh29, 8'sh0f, 8'sh01, 8'sh22, 8'sh14, 8'shff, 8'sh2a, 8'shc8, 8'shea, 8'shfd, 8'sh16
    /* (303, 0) */	    8'sh17, 8'sh17, 8'shc4, 8'shc0, 8'sh22, 8'sh2c, 8'sh10, 8'sh01, 8'sh25, 8'sh16, 8'shff, 8'sh2d, 8'shc4, 8'she8, 8'shfd, 8'sh17
    /* (304, 0) */	    8'sh18, 8'sh18, 8'shc0, 8'shbb, 8'sh25, 8'sh2f, 8'sh11, 8'sh01, 8'sh27, 8'sh17, 8'shff, 8'sh30, 8'shc0, 8'she7, 8'shfd, 8'sh19
    /* (305, 0) */	    8'sh1a, 8'sh1a, 8'shbc, 8'shb7, 8'sh27, 8'sh32, 8'sh12, 8'sh01, 8'sh29, 8'sh19, 8'shff, 8'sh33, 8'shbc, 8'she5, 8'shfc, 8'sh1a
    /* (306, 0) */	    8'sh1b, 8'sh1b, 8'shb8, 8'shb3, 8'sh29, 8'sh34, 8'sh13, 8'sh01, 8'sh2c, 8'sh1a, 8'shff, 8'sh36, 8'shb8, 8'she3, 8'shfc, 8'sh1c
    /* (307, 0) */	    8'sh1d, 8'sh1d, 8'shb4, 8'shaf, 8'sh2b, 8'sh37, 8'sh14, 8'sh01, 8'sh2e, 8'sh1c, 8'shff, 8'sh39, 8'shb4, 8'she2, 8'shfc, 8'sh1d
    /* (308, 0) */	    8'sh1f, 8'sh1f, 8'shb0, 8'shaa, 8'sh2e, 8'sh3a, 8'sh15, 8'sh01, 8'sh31, 8'sh1d, 8'shff, 8'sh3c, 8'shb0, 8'she0, 8'shfc, 8'sh1f
    /* (309, 0) */	    8'sh20, 8'sh20, 8'shac, 8'sha6, 8'sh30, 8'sh3d, 8'sh16, 8'sh01, 8'sh33, 8'sh1f, 8'shff, 8'sh3f, 8'shac, 8'shdf, 8'shfc, 8'sh20
    /* (310, 0) */	    8'sh22, 8'sh22, 8'sha8, 8'sha2, 8'sh32, 8'sh40, 8'sh17, 8'sh01, 8'sh36, 8'sh20, 8'shff, 8'sh43, 8'sha8, 8'shdd, 8'shfb, 8'sh22
    /* (311, 0) */	    8'sh23, 8'sh23, 8'sha4, 8'sh9d, 8'sh35, 8'sh43, 8'sh18, 8'sh01, 8'sh38, 8'sh22, 8'shff, 8'sh46, 8'sha4, 8'shdb, 8'shfb, 8'sh23
    /* (312, 0) */	    8'sh25, 8'sh25, 8'sha0, 8'sh99, 8'sh37, 8'sh46, 8'sh1a, 8'sh01, 8'sh3a, 8'sh23, 8'shff, 8'sh49, 8'sha0, 8'shda, 8'shfb, 8'sh25
    /* (313, 0) */	    8'sh26, 8'sh26, 8'sh9c, 8'sh95, 8'sh39, 8'sh49, 8'sh1b, 8'sh01, 8'sh3d, 8'sh24, 8'shff, 8'sh4c, 8'sh9c, 8'shd8, 8'shfb, 8'sh27
    /* (314, 0) */	    8'sh28, 8'sh28, 8'sh98, 8'sh91, 8'sh3b, 8'sh4c, 8'sh1c, 8'sh01, 8'sh3f, 8'sh26, 8'shff, 8'sh4f, 8'sh98, 8'shd7, 8'shfb, 8'sh28
    /* (315, 0) */	    8'sh29, 8'sh29, 8'sh94, 8'sh8c, 8'sh3e, 8'sh4f, 8'sh1d, 8'sh01, 8'sh42, 8'sh27, 8'shff, 8'sh52, 8'sh94, 8'shd5, 8'shfa, 8'sh2a
    /* (316, 0) */	    8'sh2b, 8'sh2b, 8'sh90, 8'sh88, 8'sh40, 8'sh52, 8'sh1e, 8'sh01, 8'sh44, 8'sh29, 8'shff, 8'sh55, 8'sh90, 8'shd3, 8'shfa, 8'sh2b
    /* (317, 0) */	    8'sh2c, 8'sh2c, 8'sh8c, 8'sh84, 8'sh42, 8'sh54, 8'sh1f, 8'sh01, 8'sh47, 8'sh2a, 8'shff, 8'sh58, 8'sh8c, 8'shd2, 8'shfa, 8'sh2d
    /* (318, 0) */	    8'sh2e, 8'sh2e, 8'sh89, 8'sh80, 8'sh45, 8'sh57, 8'sh20, 8'sh01, 8'sh49, 8'sh2c, 8'shff, 8'sh5b, 8'sh88, 8'shd0, 8'shfa, 8'sh2e
    /* (319, 0) */	    8'sh2f, 8'sh2f, 8'sh85, 8'sh80, 8'sh47, 8'sh5a, 8'sh21, 8'sh02, 8'sh4c, 8'sh2d, 8'shff, 8'sh5e, 8'sh84, 8'shcf, 8'shfa, 8'sh30
    /* (320, 0) */	    8'sh13, 8'sh80, 8'sh80, 8'sh84, 8'sh80, 8'sh80, 8'sh01, 8'sh7f, 8'sh58, 8'sh7c, 8'sh1c, 8'sh3e, 8'sh69, 8'shf7, 8'sh7f, 8'sh7f
    /* (321, 0) */	    8'sh12, 8'sh84, 8'sh84, 8'sh88, 8'sh84, 8'sh84, 8'sh01, 8'sh7c, 8'sh55, 8'sh78, 8'sh1c, 8'sh3d, 8'sh66, 8'shf8, 8'sh7c, 8'sh7c
    /* (322, 0) */	    8'sh12, 8'sh88, 8'sh88, 8'sh8c, 8'sh88, 8'sh88, 8'sh01, 8'sh78, 8'sh52, 8'sh74, 8'sh1b, 8'sh3b, 8'sh63, 8'shf8, 8'sh78, 8'sh78
    /* (323, 0) */	    8'sh11, 8'sh8c, 8'sh8c, 8'sh8f, 8'sh8c, 8'sh8c, 8'sh01, 8'sh74, 8'sh50, 8'sh70, 8'sh1a, 8'sh39, 8'sh60, 8'shf8, 8'sh74, 8'sh74
    /* (324, 0) */	    8'sh11, 8'sh90, 8'sh90, 8'sh93, 8'sh90, 8'sh90, 8'sh01, 8'sh70, 8'sh4d, 8'sh6c, 8'sh19, 8'sh37, 8'sh5c, 8'shf8, 8'sh70, 8'sh70
    /* (325, 0) */	    8'sh10, 8'sh94, 8'sh94, 8'sh97, 8'sh94, 8'sh94, 8'sh01, 8'sh6c, 8'sh4a, 8'sh68, 8'sh18, 8'sh35, 8'sh59, 8'shf9, 8'sh6c, 8'sh6c
    /* (326, 0) */	    8'sh0f, 8'sh98, 8'sh98, 8'sh9b, 8'sh98, 8'sh98, 8'sh01, 8'sh68, 8'sh47, 8'sh65, 8'sh17, 8'sh33, 8'sh56, 8'shf9, 8'sh68, 8'sh68
    /* (327, 0) */	    8'sh0f, 8'sh9c, 8'sh9c, 8'sh9f, 8'sh9c, 8'sh9c, 8'sh01, 8'sh64, 8'sh45, 8'sh61, 8'sh16, 8'sh31, 8'sh52, 8'shf9, 8'sh64, 8'sh64
    /* (328, 0) */	    8'sh0e, 8'sha0, 8'sha0, 8'sha3, 8'sha0, 8'sha0, 8'sh01, 8'sh60, 8'sh42, 8'sh5d, 8'sh15, 8'sh2f, 8'sh4f, 8'shfa, 8'sh60, 8'sh60
    /* (329, 0) */	    8'sh0e, 8'sha4, 8'sha4, 8'sha7, 8'sha4, 8'sha4, 8'sh01, 8'sh5c, 8'sh3f, 8'sh59, 8'sh14, 8'sh2d, 8'sh4c, 8'shfa, 8'sh5c, 8'sh5c
    /* (330, 0) */	    8'sh0d, 8'sha8, 8'sha8, 8'shab, 8'sha8, 8'sha8, 8'sh01, 8'sh58, 8'sh3c, 8'sh55, 8'sh14, 8'sh2b, 8'sh48, 8'shfa, 8'sh58, 8'sh58
    /* (331, 0) */	    8'sh0c, 8'shac, 8'shac, 8'shae, 8'shac, 8'shac, 8'sh01, 8'sh54, 8'sh3a, 8'sh51, 8'sh13, 8'sh29, 8'sh45, 8'shfa, 8'sh54, 8'sh54
    /* (332, 0) */	    8'sh0c, 8'shb0, 8'shb0, 8'shb2, 8'shb0, 8'shb0, 8'sh01, 8'sh50, 8'sh37, 8'sh4d, 8'sh12, 8'sh27, 8'sh42, 8'shfb, 8'sh50, 8'sh50
    /* (333, 0) */	    8'sh0b, 8'shb4, 8'shb4, 8'shb6, 8'shb4, 8'shb4, 8'sh01, 8'sh4c, 8'sh34, 8'sh49, 8'sh11, 8'sh25, 8'sh3f, 8'shfb, 8'sh4c, 8'sh4c
    /* (334, 0) */	    8'sh0b, 8'shb8, 8'shb8, 8'shba, 8'shb8, 8'shb8, 8'sh01, 8'sh48, 8'sh31, 8'sh46, 8'sh10, 8'sh23, 8'sh3b, 8'shfb, 8'sh48, 8'sh48
    /* (335, 0) */	    8'sh0a, 8'shbc, 8'shbc, 8'shbe, 8'shbc, 8'shbc, 8'sh01, 8'sh44, 8'sh2f, 8'sh42, 8'sh0f, 8'sh21, 8'sh38, 8'shfb, 8'sh44, 8'sh44
    /* (336, 0) */	    8'sh09, 8'shc0, 8'shc0, 8'shc2, 8'shc0, 8'shc0, 8'sh01, 8'sh40, 8'sh2c, 8'sh3e, 8'sh0e, 8'sh1f, 8'sh35, 8'shfc, 8'sh40, 8'sh40
    /* (337, 0) */	    8'sh09, 8'shc4, 8'shc4, 8'shc6, 8'shc4, 8'shc4, 8'sh01, 8'sh3c, 8'sh29, 8'sh3a, 8'sh0d, 8'sh1d, 8'sh31, 8'shfc, 8'sh3c, 8'sh3c
    /* (338, 0) */	    8'sh08, 8'shc8, 8'shc8, 8'shca, 8'shc8, 8'shc8, 8'sh01, 8'sh38, 8'sh26, 8'sh36, 8'sh0c, 8'sh1b, 8'sh2e, 8'shfc, 8'sh38, 8'sh38
    /* (339, 0) */	    8'sh08, 8'shcc, 8'shcc, 8'shce, 8'shcc, 8'shcc, 8'sh00, 8'sh34, 8'sh24, 8'sh32, 8'sh0c, 8'sh19, 8'sh2b, 8'shfd, 8'sh34, 8'sh34
    /* (340, 0) */	    8'sh07, 8'shd0, 8'shd0, 8'shd1, 8'shd0, 8'shd0, 8'sh00, 8'sh30, 8'sh21, 8'sh2e, 8'sh0b, 8'sh17, 8'sh28, 8'shfd, 8'sh30, 8'sh30
    /* (341, 0) */	    8'sh07, 8'shd4, 8'shd4, 8'shd5, 8'shd4, 8'shd4, 8'sh00, 8'sh2c, 8'sh1e, 8'sh2b, 8'sh0a, 8'sh15, 8'sh24, 8'shfd, 8'sh2c, 8'sh2c
    /* (342, 0) */	    8'sh06, 8'shd8, 8'shd8, 8'shd9, 8'shd8, 8'shd8, 8'sh00, 8'sh28, 8'sh1b, 8'sh27, 8'sh09, 8'sh14, 8'sh21, 8'shfd, 8'sh28, 8'sh28
    /* (343, 0) */	    8'sh05, 8'shdc, 8'shdc, 8'shdd, 8'shdc, 8'shdc, 8'sh00, 8'sh24, 8'sh19, 8'sh23, 8'sh08, 8'sh12, 8'sh1e, 8'shfe, 8'sh24, 8'sh24
    /* (344, 0) */	    8'sh05, 8'she0, 8'she0, 8'she1, 8'she0, 8'she0, 8'sh00, 8'sh20, 8'sh16, 8'sh1f, 8'sh07, 8'sh10, 8'sh1a, 8'shfe, 8'sh20, 8'sh20
    /* (345, 0) */	    8'sh04, 8'she4, 8'she4, 8'she5, 8'she4, 8'she4, 8'sh00, 8'sh1c, 8'sh13, 8'sh1b, 8'sh06, 8'sh0e, 8'sh17, 8'shfe, 8'sh1c, 8'sh1c
    /* (346, 0) */	    8'sh04, 8'she8, 8'she8, 8'she9, 8'she8, 8'she8, 8'sh00, 8'sh18, 8'sh10, 8'sh17, 8'sh05, 8'sh0c, 8'sh14, 8'shfe, 8'sh18, 8'sh18
    /* (347, 0) */	    8'sh03, 8'shec, 8'shec, 8'shed, 8'shec, 8'shec, 8'sh00, 8'sh14, 8'sh0e, 8'sh13, 8'sh04, 8'sh0a, 8'sh10, 8'shff, 8'sh14, 8'sh14
    /* (348, 0) */	    8'sh02, 8'shf0, 8'shf0, 8'shf0, 8'shf0, 8'shf0, 8'sh00, 8'sh10, 8'sh0b, 8'sh0f, 8'sh04, 8'sh08, 8'sh0d, 8'shff, 8'sh10, 8'sh10
    /* (349, 0) */	    8'sh02, 8'shf4, 8'shf4, 8'shf4, 8'shf4, 8'shf4, 8'sh00, 8'sh0c, 8'sh08, 8'sh0c, 8'sh03, 8'sh06, 8'sh0a, 8'shff, 8'sh0c, 8'sh0c
    /* (350, 0) */	    8'sh01, 8'shf8, 8'shf8, 8'shf8, 8'shf8, 8'shf8, 8'sh00, 8'sh08, 8'sh05, 8'sh08, 8'sh02, 8'sh04, 8'sh07, 8'shff, 8'sh08, 8'sh08
    /* (351, 0) */	    8'sh01, 8'shfc, 8'shfc, 8'shfc, 8'shfc, 8'shfc, 8'sh00, 8'sh04, 8'sh03, 8'sh04, 8'sh01, 8'sh02, 8'sh03, 8'sh00, 8'sh04, 8'sh04
    /* (352, 0) */	    8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00
    /* (353, 0) */	    8'shff, 8'sh04, 8'sh04, 8'sh04, 8'sh04, 8'sh04, 8'sh00, 8'shfc, 8'shfd, 8'shfc, 8'shff, 8'shfe, 8'shfd, 8'sh00, 8'shfc, 8'shfc
    /* (354, 0) */	    8'shff, 8'sh08, 8'sh08, 8'sh08, 8'sh08, 8'sh08, 8'sh00, 8'shf8, 8'shfb, 8'shf8, 8'shfe, 8'shfc, 8'shf9, 8'sh01, 8'shf8, 8'shf8
    /* (355, 0) */	    8'shfe, 8'sh0c, 8'sh0c, 8'sh0c, 8'sh0c, 8'sh0c, 8'sh00, 8'shf4, 8'shf8, 8'shf4, 8'shfd, 8'shfa, 8'shf6, 8'sh01, 8'shf4, 8'shf4
    /* (356, 0) */	    8'shfe, 8'sh10, 8'sh10, 8'sh10, 8'sh10, 8'sh10, 8'sh00, 8'shf0, 8'shf5, 8'shf1, 8'shfc, 8'shf8, 8'shf3, 8'sh01, 8'shf0, 8'shf0
    /* (357, 0) */	    8'shfd, 8'sh14, 8'sh14, 8'sh13, 8'sh14, 8'sh14, 8'sh00, 8'shec, 8'shf2, 8'shed, 8'shfc, 8'shf6, 8'shf0, 8'sh01, 8'shec, 8'shec
    /* (358, 0) */	    8'shfc, 8'sh18, 8'sh18, 8'sh17, 8'sh18, 8'sh18, 8'sh00, 8'she8, 8'shf0, 8'she9, 8'shfb, 8'shf4, 8'shec, 8'sh02, 8'she8, 8'she8
    /* (359, 0) */	    8'shfc, 8'sh1c, 8'sh1c, 8'sh1b, 8'sh1c, 8'sh1c, 8'sh00, 8'she4, 8'shed, 8'she5, 8'shfa, 8'shf2, 8'she9, 8'sh02, 8'she4, 8'she4
    /* (360, 0) */	    8'shfb, 8'sh20, 8'sh20, 8'sh1f, 8'sh20, 8'sh20, 8'sh00, 8'she0, 8'shea, 8'she1, 8'shf9, 8'shf0, 8'she6, 8'sh02, 8'she0, 8'she0
    /* (361, 0) */	    8'shfb, 8'sh24, 8'sh24, 8'sh23, 8'sh24, 8'sh24, 8'sh00, 8'shdc, 8'she7, 8'shdd, 8'shf8, 8'shee, 8'she2, 8'sh02, 8'shdc, 8'shdc
    /* (362, 0) */	    8'shfa, 8'sh28, 8'sh28, 8'sh27, 8'sh28, 8'sh28, 8'sh00, 8'shd8, 8'she5, 8'shd9, 8'shf7, 8'shec, 8'shdf, 8'sh03, 8'shd8, 8'shd8
    /* (363, 0) */	    8'shf9, 8'sh2c, 8'sh2c, 8'sh2b, 8'sh2c, 8'sh2c, 8'sh00, 8'shd4, 8'she2, 8'shd5, 8'shf6, 8'sheb, 8'shdc, 8'sh03, 8'shd4, 8'shd4
    /* (364, 0) */	    8'shf9, 8'sh30, 8'sh30, 8'sh2f, 8'sh30, 8'sh30, 8'sh00, 8'shd0, 8'shdf, 8'shd2, 8'shf5, 8'she9, 8'shd8, 8'sh03, 8'shd0, 8'shd0
    /* (365, 0) */	    8'shf8, 8'sh34, 8'sh34, 8'sh32, 8'sh34, 8'sh34, 8'sh00, 8'shcc, 8'shdc, 8'shce, 8'shf4, 8'she7, 8'shd5, 8'sh03, 8'shcc, 8'shcc
    /* (366, 0) */	    8'shf8, 8'sh38, 8'sh38, 8'sh36, 8'sh38, 8'sh38, 8'shff, 8'shc8, 8'shda, 8'shca, 8'shf4, 8'she5, 8'shd2, 8'sh04, 8'shc8, 8'shc8
    /* (367, 0) */	    8'shf7, 8'sh3c, 8'sh3c, 8'sh3a, 8'sh3c, 8'sh3c, 8'shff, 8'shc4, 8'shd7, 8'shc6, 8'shf3, 8'she3, 8'shcf, 8'sh04, 8'shc4, 8'shc4
    /* (368, 0) */	    8'shf7, 8'sh40, 8'sh40, 8'sh3e, 8'sh40, 8'sh40, 8'shff, 8'shc0, 8'shd4, 8'shc2, 8'shf2, 8'she1, 8'shcb, 8'sh04, 8'shc0, 8'shc0
    /* (369, 0) */	    8'shf6, 8'sh44, 8'sh44, 8'sh42, 8'sh44, 8'sh44, 8'shff, 8'shbc, 8'shd1, 8'shbe, 8'shf1, 8'shdf, 8'shc8, 8'sh05, 8'shbc, 8'shbc
    /* (370, 0) */	    8'shf5, 8'sh48, 8'sh48, 8'sh46, 8'sh48, 8'sh48, 8'shff, 8'shb8, 8'shcf, 8'shba, 8'shf0, 8'shdd, 8'shc5, 8'sh05, 8'shb8, 8'shb8
    /* (371, 0) */	    8'shf5, 8'sh4c, 8'sh4c, 8'sh4a, 8'sh4c, 8'sh4c, 8'shff, 8'shb4, 8'shcc, 8'shb7, 8'shef, 8'shdb, 8'shc1, 8'sh05, 8'shb4, 8'shb4
    /* (372, 0) */	    8'shf4, 8'sh50, 8'sh50, 8'sh4e, 8'sh50, 8'sh50, 8'shff, 8'shb0, 8'shc9, 8'shb3, 8'shee, 8'shd9, 8'shbe, 8'sh05, 8'shb0, 8'shb0
    /* (373, 0) */	    8'shf4, 8'sh54, 8'sh54, 8'sh52, 8'sh54, 8'sh54, 8'shff, 8'shac, 8'shc6, 8'shaf, 8'shed, 8'shd7, 8'shbb, 8'sh06, 8'shac, 8'shac
    /* (374, 0) */	    8'shf3, 8'sh58, 8'sh58, 8'sh55, 8'sh58, 8'sh58, 8'shff, 8'sha8, 8'shc4, 8'shab, 8'shec, 8'shd5, 8'shb8, 8'sh06, 8'sha8, 8'sha8
    /* (375, 0) */	    8'shf2, 8'sh5c, 8'sh5c, 8'sh59, 8'sh5c, 8'sh5c, 8'shff, 8'sha4, 8'shc1, 8'sha7, 8'shec, 8'shd3, 8'shb4, 8'sh06, 8'sha4, 8'sha4
    /* (376, 0) */	    8'shf2, 8'sh60, 8'sh60, 8'sh5d, 8'sh60, 8'sh60, 8'shff, 8'sha0, 8'shbe, 8'sha3, 8'sheb, 8'shd1, 8'shb1, 8'sh06, 8'sha0, 8'sha0
    /* (377, 0) */	    8'shf1, 8'sh64, 8'sh64, 8'sh61, 8'sh64, 8'sh64, 8'shff, 8'sh9c, 8'shbb, 8'sh9f, 8'shea, 8'shcf, 8'shae, 8'sh07, 8'sh9c, 8'sh9c
    /* (378, 0) */	    8'shf1, 8'sh68, 8'sh68, 8'sh65, 8'sh68, 8'sh68, 8'shff, 8'sh98, 8'shb9, 8'sh9b, 8'she9, 8'shcd, 8'shaa, 8'sh07, 8'sh98, 8'sh98
    /* (379, 0) */	    8'shf0, 8'sh6c, 8'sh6c, 8'sh69, 8'sh6c, 8'sh6c, 8'shff, 8'sh94, 8'shb6, 8'sh98, 8'she8, 8'shcb, 8'sha7, 8'sh07, 8'sh94, 8'sh94
    /* (380, 0) */	    8'shef, 8'sh70, 8'sh70, 8'sh6d, 8'sh70, 8'sh70, 8'shff, 8'sh90, 8'shb3, 8'sh94, 8'she7, 8'shc9, 8'sha4, 8'sh08, 8'sh90, 8'sh90
    /* (381, 0) */	    8'shef, 8'sh74, 8'sh74, 8'sh71, 8'sh74, 8'sh74, 8'shff, 8'sh8c, 8'shb0, 8'sh90, 8'she6, 8'shc7, 8'sha0, 8'sh08, 8'sh8c, 8'sh8c
    /* (382, 0) */	    8'shee, 8'sh78, 8'sh78, 8'sh74, 8'sh78, 8'sh78, 8'shff, 8'sh88, 8'shae, 8'sh8c, 8'she5, 8'shc5, 8'sh9d, 8'sh08, 8'sh88, 8'sh88
    /* (383, 0) */	    8'shee, 8'sh7c, 8'sh7c, 8'sh78, 8'sh7c, 8'sh7c, 8'shff, 8'sh84, 8'shab, 8'sh88, 8'she4, 8'shc3, 8'sh9a, 8'sh08, 8'sh84, 8'sh84
    /* (384, 0) */	    8'sh73, 8'sh03, 8'shc1, 8'sh25, 8'she7, 8'shf2, 8'shdb, 8'she8, 8'sh1b, 8'shed, 8'sh10, 8'shb7, 8'sh03, 8'sh21, 8'shde, 8'shf5
    /* (385, 0) */	    8'sh70, 8'sh03, 8'shc3, 8'sh24, 8'she8, 8'shf2, 8'shdc, 8'she9, 8'sh1a, 8'shee, 8'sh10, 8'shb9, 8'sh03, 8'sh20, 8'shdf, 8'shf5
    /* (386, 0) */	    8'sh6c, 8'sh03, 8'shc5, 8'sh23, 8'she9, 8'shf3, 8'shdd, 8'shea, 8'sh19, 8'shee, 8'sh0f, 8'shbc, 8'sh03, 8'sh1f, 8'she0, 8'shf6
    /* (387, 0) */	    8'sh69, 8'sh03, 8'shc7, 8'sh22, 8'she9, 8'shf3, 8'shde, 8'sheb, 8'sh18, 8'shef, 8'sh0f, 8'shbe, 8'sh03, 8'sh1e, 8'she1, 8'shf6
    /* (388, 0) */	    8'sh65, 8'sh03, 8'shc9, 8'sh21, 8'shea, 8'shf4, 8'she0, 8'sheb, 8'sh17, 8'shf0, 8'sh0e, 8'shc0, 8'sh03, 8'sh1d, 8'she2, 8'shf6
    /* (389, 0) */	    8'sh61, 8'sh03, 8'shcb, 8'sh20, 8'sheb, 8'shf4, 8'she1, 8'shec, 8'sh16, 8'shf0, 8'sh0e, 8'shc3, 8'sh03, 8'sh1c, 8'she3, 8'shf7
    /* (390, 0) */	    8'sh5e, 8'sh03, 8'shcd, 8'sh1e, 8'shec, 8'shf4, 8'she2, 8'shed, 8'sh16, 8'shf1, 8'sh0d, 8'shc5, 8'sh02, 8'sh1b, 8'she4, 8'shf7
    /* (391, 0) */	    8'sh5a, 8'sh03, 8'shcf, 8'sh1d, 8'shed, 8'shf5, 8'she3, 8'shee, 8'sh15, 8'shf1, 8'sh0d, 8'shc7, 8'sh02, 8'sh1a, 8'she5, 8'shf7
    /* (392, 0) */	    8'sh57, 8'sh02, 8'shd1, 8'sh1c, 8'shed, 8'shf5, 8'she4, 8'shee, 8'sh14, 8'shf2, 8'sh0c, 8'shc9, 8'sh02, 8'sh19, 8'she6, 8'shf8
    /* (393, 0) */	    8'sh53, 8'sh02, 8'shd3, 8'sh1b, 8'shee, 8'shf6, 8'she5, 8'shef, 8'sh13, 8'shf3, 8'sh0c, 8'shcc, 8'sh02, 8'sh18, 8'she7, 8'shf8
    /* (394, 0) */	    8'sh4f, 8'sh02, 8'shd5, 8'sh1a, 8'shef, 8'shf6, 8'she7, 8'shf0, 8'sh12, 8'shf3, 8'sh0b, 8'shce, 8'sh02, 8'sh17, 8'she9, 8'shf8
    /* (395, 0) */	    8'sh4c, 8'sh02, 8'shd7, 8'sh19, 8'shf0, 8'shf7, 8'she8, 8'shf1, 8'sh11, 8'shf4, 8'sh0b, 8'shd0, 8'sh02, 8'sh16, 8'shea, 8'shf9
    /* (396, 0) */	    8'sh48, 8'sh02, 8'shd9, 8'sh17, 8'shf0, 8'shf7, 8'she9, 8'shf1, 8'sh11, 8'shf4, 8'sh0a, 8'shd2, 8'sh02, 8'sh15, 8'sheb, 8'shf9
    /* (397, 0) */	    8'sh44, 8'sh02, 8'shdb, 8'sh16, 8'shf1, 8'shf8, 8'shea, 8'shf2, 8'sh10, 8'shf5, 8'sh0a, 8'shd5, 8'sh02, 8'sh14, 8'shec, 8'shf9
    /* (398, 0) */	    8'sh41, 8'sh02, 8'shdc, 8'sh15, 8'shf2, 8'shf8, 8'sheb, 8'shf3, 8'sh0f, 8'shf5, 8'sh09, 8'shd7, 8'sh02, 8'sh13, 8'shed, 8'shfa
    /* (399, 0) */	    8'sh3d, 8'sh02, 8'shde, 8'sh14, 8'shf3, 8'shf8, 8'shec, 8'shf3, 8'sh0e, 8'shf6, 8'sh09, 8'shd9, 8'sh02, 8'sh12, 8'shee, 8'shfa
    /* (400, 0) */	    8'sh3a, 8'sh02, 8'she0, 8'sh13, 8'shf4, 8'shf9, 8'shed, 8'shf4, 8'sh0d, 8'shf7, 8'sh08, 8'shdc, 8'sh01, 8'sh11, 8'shef, 8'shfb
    /* (401, 0) */	    8'sh36, 8'sh02, 8'she2, 8'sh12, 8'shf4, 8'shf9, 8'shef, 8'shf5, 8'sh0c, 8'shf7, 8'sh08, 8'shde, 8'sh01, 8'sh10, 8'shf0, 8'shfb
    /* (402, 0) */	    8'sh32, 8'sh01, 8'she4, 8'sh10, 8'shf5, 8'shfa, 8'shf0, 8'shf6, 8'sh0c, 8'shf8, 8'sh07, 8'she0, 8'sh01, 8'sh0e, 8'shf1, 8'shfb
    /* (403, 0) */	    8'sh2f, 8'sh01, 8'she6, 8'sh0f, 8'shf6, 8'shfa, 8'shf1, 8'shf6, 8'sh0b, 8'shf8, 8'sh07, 8'she2, 8'sh01, 8'sh0d, 8'shf2, 8'shfc
    /* (404, 0) */	    8'sh2b, 8'sh01, 8'she8, 8'sh0e, 8'shf7, 8'shfb, 8'shf2, 8'shf7, 8'sh0a, 8'shf9, 8'sh06, 8'she5, 8'sh01, 8'sh0c, 8'shf3, 8'shfc
    /* (405, 0) */	    8'sh28, 8'sh01, 8'shea, 8'sh0d, 8'shf7, 8'shfb, 8'shf3, 8'shf8, 8'sh09, 8'shfa, 8'sh06, 8'she7, 8'sh01, 8'sh0b, 8'shf4, 8'shfc
    /* (406, 0) */	    8'sh24, 8'sh01, 8'shec, 8'sh0c, 8'shf8, 8'shfc, 8'shf4, 8'shf9, 8'sh08, 8'shfa, 8'sh05, 8'she9, 8'sh01, 8'sh0a, 8'shf5, 8'shfd
    /* (407, 0) */	    8'sh20, 8'sh01, 8'shee, 8'sh0b, 8'shf9, 8'shfc, 8'shf6, 8'shf9, 8'sh07, 8'shfb, 8'sh05, 8'shec, 8'sh01, 8'sh09, 8'shf6, 8'shfd
    /* (408, 0) */	    8'sh1d, 8'sh01, 8'shf0, 8'sh09, 8'shfa, 8'shfc, 8'shf7, 8'shfa, 8'sh07, 8'shfb, 8'sh04, 8'shee, 8'sh01, 8'sh08, 8'shf7, 8'shfd
    /* (409, 0) */	    8'sh19, 8'sh01, 8'shf2, 8'sh08, 8'shfb, 8'shfd, 8'shf8, 8'shfb, 8'sh06, 8'shfc, 8'sh04, 8'shf0, 8'sh01, 8'sh07, 8'shf9, 8'shfe
    /* (410, 0) */	    8'sh16, 8'sh01, 8'shf4, 8'sh07, 8'shfb, 8'shfd, 8'shf9, 8'shfc, 8'sh05, 8'shfc, 8'sh03, 8'shf2, 8'sh01, 8'sh06, 8'shfa, 8'shfe
    /* (411, 0) */	    8'sh12, 8'sh01, 8'shf6, 8'sh06, 8'shfc, 8'shfe, 8'shfa, 8'shfc, 8'sh04, 8'shfd, 8'sh03, 8'shf5, 8'sh00, 8'sh05, 8'shfb, 8'shfe
    /* (412, 0) */	    8'sh0e, 8'sh00, 8'shf8, 8'sh05, 8'shfd, 8'shfe, 8'shfb, 8'shfd, 8'sh03, 8'shfe, 8'sh02, 8'shf7, 8'sh00, 8'sh04, 8'shfc, 8'shff
    /* (413, 0) */	    8'sh0b, 8'sh00, 8'shfa, 8'sh04, 8'shfe, 8'shff, 8'shfd, 8'shfe, 8'sh02, 8'shfe, 8'sh02, 8'shf9, 8'sh00, 8'sh03, 8'shfd, 8'shff
    /* (414, 0) */	    8'sh07, 8'sh00, 8'shfc, 8'sh02, 8'shfe, 8'shff, 8'shfe, 8'shff, 8'sh02, 8'shff, 8'sh01, 8'shfb, 8'sh00, 8'sh02, 8'shfe, 8'shff
    /* (415, 0) */	    8'sh04, 8'sh00, 8'shfe, 8'sh01, 8'shff, 8'sh00, 8'shff, 8'shff, 8'sh01, 8'shff, 8'sh01, 8'shfe, 8'sh00, 8'sh01, 8'shff, 8'sh00
    /* (416, 0) */	    8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00
    /* (417, 0) */	    8'shfc, 8'sh00, 8'sh02, 8'shff, 8'sh01, 8'sh00, 8'sh01, 8'sh01, 8'shff, 8'sh01, 8'shff, 8'sh02, 8'sh00, 8'shff, 8'sh01, 8'sh00
    /* (418, 0) */	    8'shf9, 8'sh00, 8'sh04, 8'shfe, 8'sh02, 8'sh01, 8'sh02, 8'sh01, 8'shfe, 8'sh01, 8'shff, 8'sh05, 8'sh00, 8'shfe, 8'sh02, 8'sh01
    /* (419, 0) */	    8'shf5, 8'sh00, 8'sh06, 8'shfc, 8'sh02, 8'sh01, 8'sh03, 8'sh02, 8'shfe, 8'sh02, 8'shfe, 8'sh07, 8'sh00, 8'shfd, 8'sh03, 8'sh01
    /* (420, 0) */	    8'shf2, 8'sh00, 8'sh08, 8'shfb, 8'sh03, 8'sh02, 8'sh05, 8'sh03, 8'shfd, 8'sh02, 8'shfe, 8'sh09, 8'sh00, 8'shfc, 8'sh04, 8'sh01
    /* (421, 0) */	    8'shee, 8'shff, 8'sh0a, 8'shfa, 8'sh04, 8'sh02, 8'sh06, 8'sh04, 8'shfc, 8'sh03, 8'shfd, 8'sh0b, 8'sh00, 8'shfb, 8'sh05, 8'sh02
    /* (422, 0) */	    8'shea, 8'shff, 8'sh0c, 8'shf9, 8'sh05, 8'sh03, 8'sh07, 8'sh04, 8'shfb, 8'sh04, 8'shfd, 8'sh0e, 8'shff, 8'shfa, 8'sh06, 8'sh02
    /* (423, 0) */	    8'she7, 8'shff, 8'sh0e, 8'shf8, 8'sh05, 8'sh03, 8'sh08, 8'sh05, 8'shfa, 8'sh04, 8'shfc, 8'sh10, 8'shff, 8'shf9, 8'sh07, 8'sh02
    /* (424, 0) */	    8'she3, 8'shff, 8'sh10, 8'shf7, 8'sh06, 8'sh04, 8'sh09, 8'sh06, 8'shf9, 8'sh05, 8'shfc, 8'sh12, 8'shff, 8'shf8, 8'sh09, 8'sh03
    /* (425, 0) */	    8'she0, 8'shff, 8'sh12, 8'shf5, 8'sh07, 8'sh04, 8'sh0a, 8'sh07, 8'shf9, 8'sh05, 8'shfb, 8'sh14, 8'shff, 8'shf7, 8'sh0a, 8'sh03
    /* (426, 0) */	    8'shdc, 8'shff, 8'sh14, 8'shf4, 8'sh08, 8'sh04, 8'sh0c, 8'sh07, 8'shf8, 8'sh06, 8'shfb, 8'sh17, 8'shff, 8'shf6, 8'sh0b, 8'sh03
    /* (427, 0) */	    8'shd8, 8'shff, 8'sh16, 8'shf3, 8'sh09, 8'sh05, 8'sh0d, 8'sh08, 8'shf7, 8'sh06, 8'shfa, 8'sh19, 8'shff, 8'shf5, 8'sh0c, 8'sh04
    /* (428, 0) */	    8'shd5, 8'shff, 8'sh18, 8'shf2, 8'sh09, 8'sh05, 8'sh0e, 8'sh09, 8'shf6, 8'sh07, 8'shfa, 8'sh1b, 8'shff, 8'shf4, 8'sh0d, 8'sh04
    /* (429, 0) */	    8'shd1, 8'shff, 8'sh1a, 8'shf1, 8'sh0a, 8'sh06, 8'sh0f, 8'sh0a, 8'shf5, 8'sh08, 8'shf9, 8'sh1e, 8'shff, 8'shf3, 8'sh0e, 8'sh04
    /* (430, 0) */	    8'shce, 8'shff, 8'sh1c, 8'shf0, 8'sh0b, 8'sh06, 8'sh10, 8'sh0a, 8'shf4, 8'sh08, 8'shf9, 8'sh20, 8'shff, 8'shf2, 8'sh0f, 8'sh05
    /* (431, 0) */	    8'shca, 8'shfe, 8'sh1e, 8'shee, 8'sh0c, 8'sh07, 8'sh11, 8'sh0b, 8'shf4, 8'sh09, 8'shf8, 8'sh22, 8'shff, 8'shf0, 8'sh10, 8'sh05
    /* (432, 0) */	    8'shc6, 8'shfe, 8'sh20, 8'shed, 8'sh0c, 8'sh07, 8'sh13, 8'sh0c, 8'shf3, 8'sh09, 8'shf8, 8'sh24, 8'shff, 8'shef, 8'sh11, 8'sh05
    /* (433, 0) */	    8'shc3, 8'shfe, 8'sh22, 8'shec, 8'sh0d, 8'sh08, 8'sh14, 8'sh0d, 8'shf2, 8'sh0a, 8'shf7, 8'sh27, 8'shfe, 8'shee, 8'sh12, 8'sh06
    /* (434, 0) */	    8'shbf, 8'shfe, 8'sh24, 8'sheb, 8'sh0e, 8'sh08, 8'sh15, 8'sh0d, 8'shf1, 8'sh0b, 8'shf7, 8'sh29, 8'shfe, 8'shed, 8'sh13, 8'sh06
    /* (435, 0) */	    8'shbc, 8'shfe, 8'sh25, 8'shea, 8'sh0f, 8'sh08, 8'sh16, 8'sh0e, 8'shf0, 8'sh0b, 8'shf6, 8'sh2b, 8'shfe, 8'shec, 8'sh14, 8'sh07
    /* (436, 0) */	    8'shb8, 8'shfe, 8'sh27, 8'she9, 8'sh10, 8'sh09, 8'sh17, 8'sh0f, 8'shef, 8'sh0c, 8'shf6, 8'sh2e, 8'shfe, 8'sheb, 8'sh15, 8'sh07
    /* (437, 0) */	    8'shb4, 8'shfe, 8'sh29, 8'she7, 8'sh10, 8'sh09, 8'sh18, 8'sh0f, 8'shef, 8'sh0c, 8'shf5, 8'sh30, 8'shfe, 8'shea, 8'sh16, 8'sh07
    /* (438, 0) */	    8'shb1, 8'shfe, 8'sh2b, 8'she6, 8'sh11, 8'sh0a, 8'sh19, 8'sh10, 8'shee, 8'sh0d, 8'shf5, 8'sh32, 8'shfe, 8'she9, 8'sh17, 8'sh08
    /* (439, 0) */	    8'shad, 8'shfe, 8'sh2d, 8'she5, 8'sh12, 8'sh0a, 8'sh1b, 8'sh11, 8'shed, 8'sh0d, 8'shf4, 8'sh34, 8'shfe, 8'she8, 8'sh19, 8'sh08
    /* (440, 0) */	    8'sha9, 8'shfe, 8'sh2f, 8'she4, 8'sh13, 8'sh0b, 8'sh1c, 8'sh12, 8'shec, 8'sh0e, 8'shf4, 8'sh37, 8'shfe, 8'she7, 8'sh1a, 8'sh08
    /* (441, 0) */	    8'sha6, 8'shfd, 8'sh31, 8'she3, 8'sh13, 8'sh0b, 8'sh1d, 8'sh12, 8'sheb, 8'sh0f, 8'shf3, 8'sh39, 8'shfe, 8'she6, 8'sh1b, 8'sh09
    /* (442, 0) */	    8'sha2, 8'shfd, 8'sh33, 8'she2, 8'sh14, 8'sh0c, 8'sh1e, 8'sh13, 8'shea, 8'sh0f, 8'shf3, 8'sh3b, 8'shfe, 8'she5, 8'sh1c, 8'sh09
    /* (443, 0) */	    8'sh9f, 8'shfd, 8'sh35, 8'she0, 8'sh15, 8'sh0c, 8'sh1f, 8'sh14, 8'shea, 8'sh10, 8'shf2, 8'sh3d, 8'shfd, 8'she4, 8'sh1d, 8'sh09
    /* (444, 0) */	    8'sh9b, 8'shfd, 8'sh37, 8'shdf, 8'sh16, 8'sh0c, 8'sh20, 8'sh15, 8'she9, 8'sh10, 8'shf2, 8'sh40, 8'shfd, 8'she3, 8'sh1e, 8'sh0a
    /* (445, 0) */	    8'sh97, 8'shfd, 8'sh39, 8'shde, 8'sh17, 8'sh0d, 8'sh22, 8'sh15, 8'she8, 8'sh11, 8'shf1, 8'sh42, 8'shfd, 8'she2, 8'sh1f, 8'sh0a
    /* (446, 0) */	    8'sh94, 8'shfd, 8'sh3b, 8'shdd, 8'sh17, 8'sh0d, 8'sh23, 8'sh16, 8'she7, 8'sh12, 8'shf1, 8'sh44, 8'shfd, 8'she1, 8'sh20, 8'sh0a
    /* (447, 0) */	    8'sh90, 8'shfd, 8'sh3d, 8'shdc, 8'sh18, 8'sh0e, 8'sh24, 8'sh17, 8'she6, 8'sh12, 8'shf0, 8'sh47, 8'shfd, 8'she0, 8'sh21, 8'sh0b
    /* (448, 0) */	    8'sh80, 8'sh42, 8'sh7f, 8'shdc, 8'sh5e, 8'sh50, 8'sh70, 8'sh29, 8'sh80, 8'sh7f, 8'sh7f, 8'sh7f, 8'sh80, 8'sh80, 8'sh7f, 8'sh31
    /* (449, 0) */	    8'sh80, 8'sh40, 8'sh7c, 8'shdd, 8'sh5c, 8'sh4d, 8'sh6d, 8'sh27, 8'sh84, 8'sh7c, 8'sh7b, 8'sh7c, 8'sh84, 8'sh84, 8'sh7b, 8'sh30
    /* (450, 0) */	    8'sh84, 8'sh3e, 8'sh78, 8'shde, 8'sh59, 8'sh4b, 8'sh69, 8'sh26, 8'sh88, 8'sh78, 8'sh77, 8'sh78, 8'sh88, 8'sh88, 8'sh77, 8'sh2e
    /* (451, 0) */	    8'sh88, 8'sh3b, 8'sh74, 8'shdf, 8'sh56, 8'sh48, 8'sh66, 8'sh25, 8'sh8c, 8'sh74, 8'sh73, 8'sh74, 8'sh8c, 8'sh8c, 8'sh74, 8'sh2d
    /* (452, 0) */	    8'sh8d, 8'sh39, 8'sh70, 8'she0, 8'sh53, 8'sh46, 8'sh62, 8'sh24, 8'sh90, 8'sh70, 8'sh70, 8'sh70, 8'sh90, 8'sh90, 8'sh70, 8'sh2b
    /* (453, 0) */	    8'sh91, 8'sh37, 8'sh6c, 8'she1, 8'sh50, 8'sh43, 8'sh5f, 8'sh22, 8'sh94, 8'sh6c, 8'sh6c, 8'sh6c, 8'sh94, 8'sh94, 8'sh6c, 8'sh29
    /* (454, 0) */	    8'sh95, 8'sh35, 8'sh68, 8'she3, 8'sh4d, 8'sh41, 8'sh5b, 8'sh21, 8'sh98, 8'sh68, 8'sh68, 8'sh68, 8'sh98, 8'sh98, 8'sh68, 8'sh28
    /* (455, 0) */	    8'sh99, 8'sh33, 8'sh64, 8'she4, 8'sh4a, 8'sh3e, 8'sh58, 8'sh20, 8'sh9c, 8'sh64, 8'sh64, 8'sh64, 8'sh9c, 8'sh9c, 8'sh64, 8'sh26
    /* (456, 0) */	    8'sh9d, 8'sh31, 8'sh60, 8'she5, 8'sh47, 8'sh3c, 8'sh54, 8'sh1e, 8'sha0, 8'sh60, 8'sh60, 8'sh60, 8'sha0, 8'sha0, 8'sh60, 8'sh25
    /* (457, 0) */	    8'sha1, 8'sh2f, 8'sh5c, 8'she6, 8'sh44, 8'sh39, 8'sh51, 8'sh1d, 8'sha4, 8'sh5c, 8'sh5c, 8'sh5c, 8'sha4, 8'sha4, 8'sh5c, 8'sh23
    /* (458, 0) */	    8'sha5, 8'sh2d, 8'sh58, 8'she7, 8'sh41, 8'sh37, 8'sh4d, 8'sh1c, 8'sha8, 8'sh58, 8'sh58, 8'sh58, 8'sha8, 8'sha8, 8'sh58, 8'sh22
    /* (459, 0) */	    8'sha9, 8'sh2b, 8'sh54, 8'she8, 8'sh3e, 8'sh34, 8'sh4a, 8'sh1b, 8'shac, 8'sh54, 8'sh54, 8'sh54, 8'shac, 8'shac, 8'sh54, 8'sh20
    /* (460, 0) */	    8'shae, 8'sh29, 8'sh50, 8'she9, 8'sh3b, 8'sh32, 8'sh46, 8'sh19, 8'shb0, 8'sh50, 8'sh50, 8'sh50, 8'shb0, 8'shb0, 8'sh50, 8'sh1f
    /* (461, 0) */	    8'shb2, 8'sh27, 8'sh4c, 8'sheb, 8'sh38, 8'sh2f, 8'sh43, 8'sh18, 8'shb4, 8'sh4c, 8'sh4c, 8'sh4c, 8'shb4, 8'shb4, 8'sh4c, 8'sh1d
    /* (462, 0) */	    8'shb6, 8'sh25, 8'sh48, 8'shec, 8'sh35, 8'sh2d, 8'sh3f, 8'sh17, 8'shb8, 8'sh48, 8'sh48, 8'sh48, 8'shb8, 8'shb8, 8'sh48, 8'sh1c
    /* (463, 0) */	    8'shba, 8'sh23, 8'sh44, 8'shed, 8'sh32, 8'sh2a, 8'sh3c, 8'sh16, 8'shbc, 8'sh44, 8'sh44, 8'sh44, 8'shbc, 8'shbc, 8'sh44, 8'sh1a
    /* (464, 0) */	    8'shbe, 8'sh21, 8'sh40, 8'shee, 8'sh2f, 8'sh28, 8'sh38, 8'sh14, 8'shc0, 8'sh40, 8'sh40, 8'sh40, 8'shc0, 8'shc0, 8'sh40, 8'sh19
    /* (465, 0) */	    8'shc2, 8'sh1f, 8'sh3c, 8'shef, 8'sh2c, 8'sh25, 8'sh35, 8'sh13, 8'shc4, 8'sh3c, 8'sh3c, 8'sh3c, 8'shc4, 8'shc4, 8'sh3c, 8'sh17
    /* (466, 0) */	    8'shc6, 8'sh1d, 8'sh38, 8'shf0, 8'sh29, 8'sh23, 8'sh31, 8'sh12, 8'shc8, 8'sh38, 8'sh38, 8'sh38, 8'shc8, 8'shc8, 8'sh38, 8'sh16
    /* (467, 0) */	    8'shca, 8'sh1b, 8'sh34, 8'shf1, 8'sh26, 8'sh20, 8'sh2e, 8'sh11, 8'shcc, 8'sh34, 8'sh34, 8'sh34, 8'shcc, 8'shcc, 8'sh34, 8'sh14
    /* (468, 0) */	    8'shcf, 8'sh19, 8'sh30, 8'shf2, 8'sh23, 8'sh1e, 8'sh2a, 8'sh0f, 8'shd0, 8'sh30, 8'sh30, 8'sh30, 8'shd0, 8'shd0, 8'sh30, 8'sh12
    /* (469, 0) */	    8'shd3, 8'sh17, 8'sh2c, 8'shf4, 8'sh20, 8'sh1b, 8'sh27, 8'sh0e, 8'shd4, 8'sh2c, 8'sh2c, 8'sh2c, 8'shd4, 8'shd4, 8'sh2c, 8'sh11
    /* (470, 0) */	    8'shd7, 8'sh15, 8'sh28, 8'shf5, 8'sh1e, 8'sh19, 8'sh23, 8'sh0d, 8'shd8, 8'sh28, 8'sh28, 8'sh28, 8'shd8, 8'shd8, 8'sh28, 8'sh0f
    /* (471, 0) */	    8'shdb, 8'sh12, 8'sh24, 8'shf6, 8'sh1b, 8'sh16, 8'sh20, 8'sh0b, 8'shdc, 8'sh24, 8'sh24, 8'sh24, 8'shdc, 8'shdc, 8'sh24, 8'sh0e
    /* (472, 0) */	    8'shdf, 8'sh10, 8'sh20, 8'shf7, 8'sh18, 8'sh14, 8'sh1c, 8'sh0a, 8'she0, 8'sh20, 8'sh20, 8'sh20, 8'she0, 8'she0, 8'sh20, 8'sh0c
    /* (473, 0) */	    8'she3, 8'sh0e, 8'sh1c, 8'shf8, 8'sh15, 8'sh11, 8'sh19, 8'sh09, 8'she4, 8'sh1c, 8'sh1c, 8'sh1c, 8'she4, 8'she4, 8'sh1c, 8'sh0b
    /* (474, 0) */	    8'she7, 8'sh0c, 8'sh18, 8'shf9, 8'sh12, 8'sh0f, 8'sh15, 8'sh08, 8'she8, 8'sh18, 8'sh18, 8'sh18, 8'she8, 8'she8, 8'sh18, 8'sh09
    /* (475, 0) */	    8'sheb, 8'sh0a, 8'sh14, 8'shfa, 8'sh0f, 8'sh0c, 8'sh12, 8'sh06, 8'shec, 8'sh14, 8'sh14, 8'sh14, 8'shec, 8'shec, 8'sh14, 8'sh08
    /* (476, 0) */	    8'shf0, 8'sh08, 8'sh10, 8'shfb, 8'sh0c, 8'sh0a, 8'sh0e, 8'sh05, 8'shf0, 8'sh10, 8'sh10, 8'sh10, 8'shf0, 8'shf0, 8'sh10, 8'sh06
    /* (477, 0) */	    8'shf4, 8'sh06, 8'sh0c, 8'shfd, 8'sh09, 8'sh07, 8'sh0b, 8'sh04, 8'shf4, 8'sh0c, 8'sh0c, 8'sh0c, 8'shf4, 8'shf4, 8'sh0c, 8'sh05
    /* (478, 0) */	    8'shf8, 8'sh04, 8'sh08, 8'shfe, 8'sh06, 8'sh05, 8'sh07, 8'sh03, 8'shf8, 8'sh08, 8'sh08, 8'sh08, 8'shf8, 8'shf8, 8'sh08, 8'sh03
    /* (479, 0) */	    8'shfc, 8'sh02, 8'sh04, 8'shff, 8'sh03, 8'sh02, 8'sh04, 8'sh01, 8'shfc, 8'sh04, 8'sh04, 8'sh04, 8'shfc, 8'shfc, 8'sh04, 8'sh02
    /* (480, 0) */	    8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00
    /* (481, 0) */	    8'sh04, 8'shfe, 8'shfc, 8'sh01, 8'shfd, 8'shfe, 8'shfc, 8'shff, 8'sh04, 8'shfc, 8'shfc, 8'shfc, 8'sh04, 8'sh04, 8'shfc, 8'shfe
    /* (482, 0) */	    8'sh08, 8'shfc, 8'shf8, 8'sh02, 8'shfa, 8'shfb, 8'shf9, 8'shfd, 8'sh08, 8'shf8, 8'shf8, 8'shf8, 8'sh08, 8'sh08, 8'shf8, 8'shfd
    /* (483, 0) */	    8'sh0c, 8'shfa, 8'shf4, 8'sh03, 8'shf7, 8'shf9, 8'shf5, 8'shfc, 8'sh0c, 8'shf4, 8'shf4, 8'shf4, 8'sh0c, 8'sh0c, 8'shf4, 8'shfb
    /* (484, 0) */	    8'sh10, 8'shf8, 8'shf0, 8'sh05, 8'shf4, 8'shf6, 8'shf2, 8'shfb, 8'sh10, 8'shf0, 8'shf0, 8'shf0, 8'sh10, 8'sh10, 8'shf0, 8'shfa
    /* (485, 0) */	    8'sh15, 8'shf6, 8'shec, 8'sh06, 8'shf1, 8'shf4, 8'shee, 8'shfa, 8'sh14, 8'shec, 8'shec, 8'shec, 8'sh14, 8'sh14, 8'shec, 8'shf8
    /* (486, 0) */	    8'sh19, 8'shf4, 8'she8, 8'sh07, 8'shee, 8'shf1, 8'sheb, 8'shf8, 8'sh18, 8'she8, 8'she8, 8'she8, 8'sh18, 8'sh18, 8'she8, 8'shf7
    /* (487, 0) */	    8'sh1d, 8'shf2, 8'she4, 8'sh08, 8'sheb, 8'shef, 8'she7, 8'shf7, 8'sh1c, 8'she4, 8'she4, 8'she4, 8'sh1c, 8'sh1c, 8'she4, 8'shf5
    /* (488, 0) */	    8'sh21, 8'shf0, 8'she0, 8'sh09, 8'she8, 8'shec, 8'she4, 8'shf6, 8'sh20, 8'she0, 8'she0, 8'she0, 8'sh20, 8'sh20, 8'she0, 8'shf4
    /* (489, 0) */	    8'sh25, 8'shee, 8'shdc, 8'sh0a, 8'she5, 8'shea, 8'she0, 8'shf5, 8'sh24, 8'shdc, 8'shdc, 8'shdc, 8'sh24, 8'sh24, 8'shdc, 8'shf2
    /* (490, 0) */	    8'sh29, 8'sheb, 8'shd8, 8'sh0b, 8'she2, 8'she7, 8'shdd, 8'shf3, 8'sh28, 8'shd8, 8'shd8, 8'shd8, 8'sh28, 8'sh28, 8'shd8, 8'shf1
    /* (491, 0) */	    8'sh2d, 8'she9, 8'shd4, 8'sh0c, 8'she0, 8'she5, 8'shd9, 8'shf2, 8'sh2c, 8'shd4, 8'shd4, 8'shd4, 8'sh2c, 8'sh2c, 8'shd4, 8'shef
    /* (492, 0) */	    8'sh31, 8'she7, 8'shd0, 8'sh0e, 8'shdd, 8'she2, 8'shd6, 8'shf1, 8'sh30, 8'shd0, 8'shd0, 8'shd0, 8'sh30, 8'sh30, 8'shd0, 8'shee
    /* (493, 0) */	    8'sh36, 8'she5, 8'shcc, 8'sh0f, 8'shda, 8'she0, 8'shd2, 8'shef, 8'sh34, 8'shcc, 8'shcc, 8'shcc, 8'sh34, 8'sh34, 8'shcc, 8'shec
    /* (494, 0) */	    8'sh3a, 8'she3, 8'shc8, 8'sh10, 8'shd7, 8'shdd, 8'shcf, 8'shee, 8'sh38, 8'shc8, 8'shc8, 8'shc8, 8'sh38, 8'sh38, 8'shc8, 8'shea
    /* (495, 0) */	    8'sh3e, 8'she1, 8'shc4, 8'sh11, 8'shd4, 8'shdb, 8'shcb, 8'shed, 8'sh3c, 8'shc4, 8'shc4, 8'shc4, 8'sh3c, 8'sh3c, 8'shc4, 8'she9
    /* (496, 0) */	    8'sh42, 8'shdf, 8'shc0, 8'sh12, 8'shd1, 8'shd8, 8'shc8, 8'shec, 8'sh40, 8'shc0, 8'shc0, 8'shc0, 8'sh40, 8'sh40, 8'shc0, 8'she7
    /* (497, 0) */	    8'sh46, 8'shdd, 8'shbc, 8'sh13, 8'shce, 8'shd6, 8'shc4, 8'shea, 8'sh44, 8'shbc, 8'shbc, 8'shbc, 8'sh44, 8'sh44, 8'shbc, 8'she6
    /* (498, 0) */	    8'sh4a, 8'shdb, 8'shb8, 8'sh14, 8'shcb, 8'shd3, 8'shc1, 8'she9, 8'sh48, 8'shb8, 8'shb8, 8'shb8, 8'sh48, 8'sh48, 8'shb8, 8'she4
    /* (499, 0) */	    8'sh4e, 8'shd9, 8'shb4, 8'sh15, 8'shc8, 8'shd1, 8'shbd, 8'she8, 8'sh4c, 8'shb4, 8'shb4, 8'shb4, 8'sh4c, 8'sh4c, 8'shb4, 8'she3
    /* (500, 0) */	    8'sh52, 8'shd7, 8'shb0, 8'sh17, 8'shc5, 8'shce, 8'shba, 8'she7, 8'sh50, 8'shb0, 8'shb0, 8'shb0, 8'sh50, 8'sh50, 8'shb0, 8'she1
    /* (501, 0) */	    8'sh57, 8'shd5, 8'shac, 8'sh18, 8'shc2, 8'shcc, 8'shb6, 8'she5, 8'sh54, 8'shac, 8'shac, 8'shac, 8'sh54, 8'sh54, 8'shac, 8'she0
    /* (502, 0) */	    8'sh5b, 8'shd3, 8'sha8, 8'sh19, 8'shbf, 8'shc9, 8'shb3, 8'she4, 8'sh58, 8'sha8, 8'sha8, 8'sha8, 8'sh58, 8'sh58, 8'sha8, 8'shde
    /* (503, 0) */	    8'sh5f, 8'shd1, 8'sha4, 8'sh1a, 8'shbc, 8'shc7, 8'shaf, 8'she3, 8'sh5c, 8'sha4, 8'sha4, 8'sha4, 8'sh5c, 8'sh5c, 8'sha4, 8'shdd
    /* (504, 0) */	    8'sh63, 8'shcf, 8'sha0, 8'sh1b, 8'shb9, 8'shc4, 8'shac, 8'she2, 8'sh60, 8'sha0, 8'sha0, 8'sha0, 8'sh60, 8'sh60, 8'sha0, 8'shdb
    /* (505, 0) */	    8'sh67, 8'shcd, 8'sh9c, 8'sh1c, 8'shb6, 8'shc2, 8'sha8, 8'she0, 8'sh64, 8'sh9c, 8'sh9c, 8'sh9c, 8'sh64, 8'sh64, 8'sh9c, 8'shda
    /* (506, 0) */	    8'sh6b, 8'shcb, 8'sh98, 8'sh1d, 8'shb3, 8'shbf, 8'sha5, 8'shdf, 8'sh68, 8'sh98, 8'sh98, 8'sh98, 8'sh68, 8'sh68, 8'sh98, 8'shd8
    /* (507, 0) */	    8'sh6f, 8'shc9, 8'sh94, 8'sh1f, 8'shb0, 8'shbd, 8'sha1, 8'shde, 8'sh6c, 8'sh94, 8'sh94, 8'sh94, 8'sh6c, 8'sh6c, 8'sh94, 8'shd7
    /* (508, 0) */	    8'sh73, 8'shc7, 8'sh90, 8'sh20, 8'shad, 8'shba, 8'sh9e, 8'shdc, 8'sh70, 8'sh90, 8'sh90, 8'sh90, 8'sh70, 8'sh70, 8'sh90, 8'shd5
    /* (509, 0) */	    8'sh78, 8'shc5, 8'sh8c, 8'sh21, 8'shaa, 8'shb8, 8'sh9a, 8'shdb, 8'sh74, 8'sh8c, 8'sh8d, 8'sh8c, 8'sh74, 8'sh74, 8'sh8c, 8'shd3
    /* (510, 0) */	    8'sh7c, 8'shc2, 8'sh88, 8'sh22, 8'sha7, 8'shb5, 8'sh97, 8'shda, 8'sh78, 8'sh88, 8'sh89, 8'sh88, 8'sh78, 8'sh78, 8'sh89, 8'shd2
    /* (511, 0) */	    8'sh7f, 8'shc0, 8'sh84, 8'sh23, 8'sha4, 8'shb3, 8'sh93, 8'shd9, 8'sh7c, 8'sh84, 8'sh85, 8'sh84, 8'sh7c, 8'sh7c, 8'sh85, 8'shd0
    /* (512, 0) */	    8'sh7f, 8'sh4f, 8'sh35, 8'sh7f, 8'sh7f, 8'sh7f, 8'sh7f, 8'sh4e, 8'sh7f, 8'shc5, 8'sh7b, 8'sh17, 8'sh7f, 8'sh2e, 8'sh7f, 8'sh7c
    /* (513, 0) */	    8'sh7f, 8'sh4d, 8'sh34, 8'sh7f, 8'sh7f, 8'sh7f, 8'sh7f, 8'sh4b, 8'sh7f, 8'shc6, 8'sh77, 8'sh17, 8'sh7f, 8'sh2c, 8'sh7f, 8'sh79
    /* (514, 0) */	    8'sh7f, 8'sh4b, 8'sh32, 8'sh7f, 8'sh7f, 8'sh7f, 8'sh7f, 8'sh49, 8'sh7f, 8'shc8, 8'sh73, 8'sh16, 8'sh7f, 8'sh2b, 8'sh7f, 8'sh75
    /* (515, 0) */	    8'sh7f, 8'sh48, 8'sh30, 8'sh7f, 8'sh7f, 8'sh7f, 8'sh7c, 8'sh46, 8'sh7c, 8'shca, 8'sh6f, 8'sh15, 8'sh7d, 8'sh2a, 8'sh7f, 8'sh71
    /* (516, 0) */	    8'sh7f, 8'sh46, 8'sh2f, 8'sh7f, 8'sh7f, 8'sh7f, 8'sh78, 8'sh44, 8'sh78, 8'shcc, 8'sh6c, 8'sh15, 8'sh79, 8'sh28, 8'sh7f, 8'sh6d
    /* (517, 0) */	    8'sh7f, 8'sh43, 8'sh2d, 8'sh7f, 8'sh7f, 8'sh7f, 8'sh73, 8'sh42, 8'sh74, 8'shce, 8'sh68, 8'sh14, 8'sh75, 8'sh27, 8'sh7f, 8'sh69
    /* (518, 0) */	    8'sh7f, 8'sh41, 8'sh2b, 8'sh7f, 8'sh7f, 8'sh7f, 8'sh6f, 8'sh3f, 8'sh6f, 8'shd0, 8'sh64, 8'sh13, 8'sh70, 8'sh25, 8'sh7f, 8'sh65
    /* (519, 0) */	    8'sh7f, 8'sh3e, 8'sh2a, 8'sh7f, 8'sh7f, 8'sh7f, 8'sh6b, 8'sh3d, 8'sh6b, 8'shd2, 8'sh60, 8'sh12, 8'sh6c, 8'sh24, 8'sh7f, 8'sh61
    /* (520, 0) */	    8'sh7f, 8'sh3c, 8'sh28, 8'sh7f, 8'sh7f, 8'sh7f, 8'sh67, 8'sh3a, 8'sh67, 8'shd3, 8'sh5c, 8'sh12, 8'sh68, 8'sh22, 8'sh7d, 8'sh5d
    /* (521, 0) */	    8'sh7f, 8'sh39, 8'sh26, 8'sh7f, 8'sh7f, 8'sh7f, 8'sh62, 8'sh38, 8'sh63, 8'shd5, 8'sh58, 8'sh11, 8'sh63, 8'sh21, 8'sh78, 8'sh59
    /* (522, 0) */	    8'sh7f, 8'sh37, 8'sh25, 8'sh7f, 8'sh7d, 8'sh7f, 8'sh5e, 8'sh35, 8'sh5e, 8'shd7, 8'sh55, 8'sh10, 8'sh5f, 8'sh20, 8'sh73, 8'sh56
    /* (523, 0) */	    8'sh7f, 8'sh34, 8'sh23, 8'sh7f, 8'sh77, 8'sh7f, 8'sh5a, 8'sh33, 8'sh5a, 8'shd9, 8'sh51, 8'sh0f, 8'sh5b, 8'sh1e, 8'sh6d, 8'sh52
    /* (524, 0) */	    8'sh7f, 8'sh32, 8'sh21, 8'sh7f, 8'sh71, 8'sh7f, 8'sh55, 8'sh31, 8'sh56, 8'shdb, 8'sh4d, 8'sh0f, 8'sh56, 8'sh1d, 8'sh68, 8'sh4e
    /* (525, 0) */	    8'sh7f, 8'sh2f, 8'sh20, 8'sh7f, 8'sh6c, 8'sh7f, 8'sh51, 8'sh2e, 8'sh51, 8'shdd, 8'sh49, 8'sh0e, 8'sh52, 8'sh1b, 8'sh63, 8'sh4a
    /* (526, 0) */	    8'sh7f, 8'sh2d, 8'sh1e, 8'sh7f, 8'sh66, 8'sh7c, 8'sh4d, 8'sh2c, 8'sh4d, 8'shdf, 8'sh45, 8'sh0d, 8'sh4e, 8'sh1a, 8'sh5e, 8'sh46
    /* (527, 0) */	    8'sh7f, 8'sh2a, 8'sh1c, 8'sh78, 8'sh60, 8'sh75, 8'sh49, 8'sh29, 8'sh49, 8'she0, 8'sh41, 8'sh0c, 8'sh49, 8'sh18, 8'sh59, 8'sh42
    /* (528, 0) */	    8'sh7f, 8'sh28, 8'sh1b, 8'sh71, 8'sh5b, 8'sh6e, 8'sh44, 8'sh27, 8'sh45, 8'she2, 8'sh3d, 8'sh0c, 8'sh45, 8'sh17, 8'sh53, 8'sh3e
    /* (529, 0) */	    8'sh7f, 8'sh25, 8'sh19, 8'sh6a, 8'sh55, 8'sh67, 8'sh40, 8'sh24, 8'sh40, 8'she4, 8'sh3a, 8'sh0b, 8'sh41, 8'sh15, 8'sh4e, 8'sh3a
    /* (530, 0) */	    8'sh7c, 8'sh23, 8'sh17, 8'sh63, 8'sh4f, 8'sh60, 8'sh3c, 8'sh22, 8'sh3c, 8'she6, 8'sh36, 8'sh0a, 8'sh3c, 8'sh14, 8'sh49, 8'sh36
    /* (531, 0) */	    8'sh73, 8'sh20, 8'sh16, 8'sh5c, 8'sh4a, 8'sh59, 8'sh38, 8'sh20, 8'sh38, 8'she8, 8'sh32, 8'sh0a, 8'sh38, 8'sh13, 8'sh44, 8'sh33
    /* (532, 0) */	    8'sh6a, 8'sh1e, 8'sh14, 8'sh55, 8'sh44, 8'sh52, 8'sh33, 8'sh1d, 8'sh33, 8'shea, 8'sh2e, 8'sh09, 8'sh34, 8'sh11, 8'sh3e, 8'sh2f
    /* (533, 0) */	    8'sh61, 8'sh1b, 8'sh12, 8'sh4e, 8'sh3e, 8'sh4c, 8'sh2f, 8'sh1b, 8'sh2f, 8'shec, 8'sh2a, 8'sh08, 8'sh2f, 8'sh10, 8'sh39, 8'sh2b
    /* (534, 0) */	    8'sh58, 8'sh19, 8'sh11, 8'sh47, 8'sh39, 8'sh45, 8'sh2b, 8'sh18, 8'sh2b, 8'shed, 8'sh26, 8'sh07, 8'sh2b, 8'sh0e, 8'sh34, 8'sh27
    /* (535, 0) */	    8'sh4f, 8'sh16, 8'sh0f, 8'sh3f, 8'sh33, 8'sh3e, 8'sh26, 8'sh16, 8'sh27, 8'shef, 8'sh23, 8'sh07, 8'sh27, 8'sh0d, 8'sh2f, 8'sh23
    /* (536, 0) */	    8'sh47, 8'sh14, 8'sh0d, 8'sh38, 8'sh2d, 8'sh37, 8'sh22, 8'sh13, 8'sh22, 8'shf1, 8'sh1f, 8'sh06, 8'sh23, 8'sh0b, 8'sh2a, 8'sh1f
    /* (537, 0) */	    8'sh3e, 8'sh11, 8'sh0c, 8'sh31, 8'sh28, 8'sh30, 8'sh1e, 8'sh11, 8'sh1e, 8'shf3, 8'sh1b, 8'sh05, 8'sh1e, 8'sh0a, 8'sh24, 8'sh1b
    /* (538, 0) */	    8'sh35, 8'sh0f, 8'sh0a, 8'sh2a, 8'sh22, 8'sh29, 8'sh1a, 8'sh0f, 8'sh1a, 8'shf5, 8'sh17, 8'sh04, 8'sh1a, 8'sh09, 8'sh1f, 8'sh17
    /* (539, 0) */	    8'sh2c, 8'sh0c, 8'sh08, 8'sh23, 8'sh1c, 8'sh22, 8'sh15, 8'sh0c, 8'sh15, 8'shf7, 8'sh13, 8'sh04, 8'sh16, 8'sh07, 8'sh1a, 8'sh13
    /* (540, 0) */	    8'sh23, 8'sh0a, 8'sh07, 8'sh1c, 8'sh17, 8'sh1b, 8'sh11, 8'sh0a, 8'sh11, 8'shf9, 8'sh0f, 8'sh03, 8'sh11, 8'sh06, 8'sh15, 8'sh10
    /* (541, 0) */	    8'sh1a, 8'sh07, 8'sh05, 8'sh15, 8'sh11, 8'sh15, 8'sh0d, 8'sh07, 8'sh0d, 8'shfa, 8'sh0c, 8'sh02, 8'sh0d, 8'sh04, 8'sh10, 8'sh0c
    /* (542, 0) */	    8'sh12, 8'sh05, 8'sh03, 8'sh0e, 8'sh0b, 8'sh0e, 8'sh09, 8'sh05, 8'sh09, 8'shfc, 8'sh08, 8'sh01, 8'sh09, 8'sh03, 8'sh0a, 8'sh08
    /* (543, 0) */	    8'sh09, 8'sh02, 8'sh02, 8'sh07, 8'sh06, 8'sh07, 8'sh04, 8'sh02, 8'sh04, 8'shfe, 8'sh04, 8'sh01, 8'sh04, 8'sh01, 8'sh05, 8'sh04
    /* (544, 0) */	    8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00, 8'sh00
    /* (545, 0) */	    8'shf7, 8'shfe, 8'shfe, 8'shf9, 8'shfa, 8'shf9, 8'shfc, 8'shfe, 8'shfc, 8'sh02, 8'shfc, 8'shff, 8'shfc, 8'shff, 8'shfb, 8'shfc
    /* (546, 0) */	    8'shee, 8'shfb, 8'shfd, 8'shf2, 8'shf5, 8'shf2, 8'shf7, 8'shfb, 8'shf7, 8'sh04, 8'shf8, 8'shff, 8'shf7, 8'shfd, 8'shf6, 8'shf8
    /* (547, 0) */	    8'she6, 8'shf9, 8'shfb, 8'sheb, 8'shef, 8'sheb, 8'shf3, 8'shf9, 8'shf3, 8'sh06, 8'shf4, 8'shfe, 8'shf3, 8'shfc, 8'shf0, 8'shf4
    /* (548, 0) */	    8'shdd, 8'shf6, 8'shf9, 8'she4, 8'she9, 8'she5, 8'shef, 8'shf6, 8'shef, 8'sh07, 8'shf1, 8'shfd, 8'shef, 8'shfa, 8'sheb, 8'shf0
    /* (549, 0) */	    8'shd4, 8'shf4, 8'shf8, 8'shdd, 8'she4, 8'shde, 8'sheb, 8'shf4, 8'sheb, 8'sh09, 8'shed, 8'shfc, 8'shea, 8'shf9, 8'she6, 8'shed
    /* (550, 0) */	    8'shcb, 8'shf1, 8'shf6, 8'shd6, 8'shde, 8'shd7, 8'she6, 8'shf1, 8'she6, 8'sh0b, 8'she9, 8'shfc, 8'she6, 8'shf7, 8'she1, 8'she9
    /* (551, 0) */	    8'shc2, 8'shef, 8'shf4, 8'shcf, 8'shd8, 8'shd0, 8'she2, 8'shef, 8'she2, 8'sh0d, 8'she5, 8'shfb, 8'she2, 8'shf6, 8'shdc, 8'she5
    /* (552, 0) */	    8'shb9, 8'shec, 8'shf3, 8'shc8, 8'shd3, 8'shc9, 8'shde, 8'shed, 8'shde, 8'sh0f, 8'she1, 8'shfa, 8'shdd, 8'shf5, 8'shd6, 8'she1
    /* (553, 0) */	    8'shb1, 8'shea, 8'shf1, 8'shc1, 8'shcd, 8'shc2, 8'shda, 8'shea, 8'shd9, 8'sh11, 8'shdd, 8'shf9, 8'shd9, 8'shf3, 8'shd1, 8'shdd
    /* (554, 0) */	    8'sha8, 8'she7, 8'shef, 8'shb9, 8'shc7, 8'shbb, 8'shd5, 8'she8, 8'shd5, 8'sh13, 8'shda, 8'shf9, 8'shd5, 8'shf2, 8'shcc, 8'shd9
    /* (555, 0) */	    8'sh9f, 8'she5, 8'shee, 8'shb2, 8'shc2, 8'shb4, 8'shd1, 8'she5, 8'shd1, 8'sh14, 8'shd6, 8'shf8, 8'shd1, 8'shf0, 8'shc7, 8'shd5
    /* (556, 0) */	    8'sh96, 8'she2, 8'shec, 8'shab, 8'shbc, 8'shae, 8'shcd, 8'she3, 8'shcd, 8'sh16, 8'shd2, 8'shf7, 8'shcc, 8'shef, 8'shc2, 8'shd1
    /* (557, 0) */	    8'sh8d, 8'she0, 8'shea, 8'sha4, 8'shb6, 8'sha7, 8'shc8, 8'she0, 8'shc8, 8'sh18, 8'shce, 8'shf6, 8'shc8, 8'shed, 8'shbc, 8'shcd
    /* (558, 0) */	    8'sh84, 8'shdd, 8'she9, 8'sh9d, 8'shb1, 8'sha0, 8'shc4, 8'shde, 8'shc4, 8'sh1a, 8'shca, 8'shf6, 8'shc4, 8'shec, 8'shb7, 8'shca
    /* (559, 0) */	    8'sh80, 8'shdb, 8'she7, 8'sh96, 8'shab, 8'sh99, 8'shc0, 8'shdc, 8'shc0, 8'sh1c, 8'shc6, 8'shf5, 8'shbf, 8'sheb, 8'shb2, 8'shc6
    /* (560, 0) */	    8'sh80, 8'shd8, 8'she5, 8'sh8f, 8'sha5, 8'sh92, 8'shbc, 8'shd9, 8'shbb, 8'sh1e, 8'shc3, 8'shf4, 8'shbb, 8'she9, 8'shad, 8'shc2
    /* (561, 0) */	    8'sh80, 8'shd6, 8'she4, 8'sh88, 8'sha0, 8'sh8b, 8'shb7, 8'shd7, 8'shb7, 8'sh20, 8'shbf, 8'shf4, 8'shb7, 8'she8, 8'sha7, 8'shbe
    /* (562, 0) */	    8'sh80, 8'shd3, 8'she2, 8'sh81, 8'sh9a, 8'sh84, 8'shb3, 8'shd4, 8'shb3, 8'sh21, 8'shbb, 8'shf3, 8'shb2, 8'she6, 8'sha2, 8'shba
    /* (563, 0) */	    8'sh80, 8'shd1, 8'she0, 8'sh80, 8'sh94, 8'sh80, 8'shaf, 8'shd2, 8'shaf, 8'sh23, 8'shb7, 8'shf2, 8'shae, 8'she5, 8'sh9d, 8'shb6
    /* (564, 0) */	    8'sh80, 8'shce, 8'shdf, 8'sh80, 8'sh8f, 8'sh80, 8'shab, 8'shcf, 8'shaa, 8'sh25, 8'shb3, 8'shf1, 8'shaa, 8'she3, 8'sh98, 8'shb2
    /* (565, 0) */	    8'sh80, 8'shcc, 8'shdd, 8'sh80, 8'sh89, 8'sh80, 8'sha6, 8'shcd, 8'sha6, 8'sh27, 8'shaf, 8'shf1, 8'sha5, 8'she2, 8'sh93, 8'shae
    /* (566, 0) */	    8'sh80, 8'shc9, 8'shdb, 8'sh80, 8'sh83, 8'sh80, 8'sha2, 8'shcb, 8'sha2, 8'sh29, 8'shab, 8'shf0, 8'sha1, 8'she0, 8'sh8d, 8'shaa
    /* (567, 0) */	    8'sh80, 8'shc7, 8'shda, 8'sh80, 8'sh80, 8'sh80, 8'sh9e, 8'shc8, 8'sh9d, 8'sh2b, 8'sha8, 8'shef, 8'sh9d, 8'shdf, 8'sh88, 8'sha7
    /* (568, 0) */	    8'sh80, 8'shc4, 8'shd8, 8'sh80, 8'sh80, 8'sh80, 8'sh99, 8'shc6, 8'sh99, 8'sh2d, 8'sha4, 8'shee, 8'sh98, 8'shde, 8'sh83, 8'sha3
    /* (569, 0) */	    8'sh80, 8'shc2, 8'shd6, 8'sh80, 8'sh80, 8'sh80, 8'sh95, 8'shc3, 8'sh95, 8'sh2e, 8'sha0, 8'shee, 8'sh94, 8'shdc, 8'sh80, 8'sh9f
    /* (570, 0) */	    8'sh80, 8'shbf, 8'shd5, 8'sh80, 8'sh80, 8'sh80, 8'sh91, 8'shc1, 8'sh91, 8'sh30, 8'sh9c, 8'shed, 8'sh90, 8'shdb, 8'sh80, 8'sh9b
    /* (571, 0) */	    8'sh80, 8'shbd, 8'shd3, 8'sh80, 8'sh80, 8'sh80, 8'sh8d, 8'shbe, 8'sh8c, 8'sh32, 8'sh98, 8'shec, 8'sh8b, 8'shd9, 8'sh80, 8'sh97
    /* (572, 0) */	    8'sh80, 8'shba, 8'shd1, 8'sh80, 8'sh80, 8'sh80, 8'sh88, 8'shbc, 8'sh88, 8'sh34, 8'sh94, 8'sheb, 8'sh87, 8'shd8, 8'sh80, 8'sh93
    /* (573, 0) */	    8'sh80, 8'shb8, 8'shd0, 8'sh80, 8'sh80, 8'sh80, 8'sh84, 8'shba, 8'sh84, 8'sh36, 8'sh91, 8'sheb, 8'sh83, 8'shd6, 8'sh80, 8'sh8f
    /* (574, 0) */	    8'sh80, 8'shb5, 8'shce, 8'sh80, 8'sh80, 8'sh80, 8'sh80, 8'shb7, 8'sh80, 8'sh38, 8'sh8d, 8'shea, 8'sh80, 8'shd5, 8'sh80, 8'sh8b
    /* (575, 0) */	    8'sh80, 8'shb3, 8'shcc, 8'sh80, 8'sh80, 8'sh80, 8'sh80, 8'shb5, 8'sh80, 8'sh3a, 8'sh89, 8'she9, 8'sh80, 8'shd4, 8'sh80, 8'sh87
};

    // 批量读取控制逻辑（优化版）
    typedef enum logic {IDLE, ACTIVE} burst_state_t;
    burst_state_t state;

    logic [4:0] counter;  // 增加1bit防止溢出

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= IDLE;
            counter <= 0;
            burst_done <= 0;
        end else begin
            case (state)
                IDLE: begin
                    burst_done <= 0;
                    if (burst_start) begin
                        state <= ACTIVE;
                        counter <= 16;  // 递减计数器
                    end
                end
                
                ACTIVE: begin
                    counter <= counter - 1;
                    if (counter == 1) begin
                        state <= IDLE;
                        burst_done <= 1;
                    end
                end
            endcase
        end
    end

    // 并行读取流水线（优化时序）
    logic [13:0] addr_reg [0:15];

    generate
        for (genvar i = 0; i < 16; i++) begin : pipeline
            // 地址计算级
            always_ff @(posedge clk) begin
                if (state == IDLE && burst_start) begin
                    addr_reg[i] <= base_addr + i;
                end else if (state == ACTIVE) begin
                    addr_reg[i] <= addr_reg[i] + 16;
                end
            end
            
            // 数据输出级
            always_ff @(posedge clk) begin
                data[i] <= lut_mem[addr_reg[i]];
            end
        end
    endgenerate

endmodule

