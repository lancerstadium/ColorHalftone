/**
 * Module       : LUTTable
 * Input        : x[31:0] - Signed/Unsigned 8-bit interger
 * Output       : y[31:0] - Unsigned/Signed 8-bit interger
 * Description  : LUT Table for read and write.
 * Author       : lancerstadium
 * Date         : Tue Mar  4 16:41:09 CST 2025
 * License      : MIT
 */

module LUTTable_x4_4b_i8_s1_D_H6 (
    input  logic        en_write,                           // 脉冲启动批量写入
    input  logic        en_read,                            // 脉冲启动批量读取
    input  logic        [9:0] base,    // 非展平基地址
    input  logic        [31:0] wdata [0:3],    // 并行输入
    output logic        [31:0] rdata [0:3]     // 并行输出
);

    // Original Shape <int8x4>: (576, 4), Total Entries: 576
    logic [31:0] lut_mem [0:2303]
    =
    '{
    /* (0, 0) */	    32'hE1190BFB, 32'hFEE7F311, 32'hFD07EA03, 32'hFE1AFD0E, 
    /* (1, 0) */	    32'hE2180BFC, 32'hFEE7F410, 32'hFD07EB03, 32'hFE19FD0E, 
    /* (2, 0) */	    32'hE3180AFC, 32'hFEE8F410, 32'hFD07EC03, 32'hFE18FE0E, 
    /* (3, 0) */	    32'hE4170AFC, 32'hFEE9F50F, 32'hFE07EC03, 32'hFF17FE0D, 
    /* (4, 0) */	    32'hE51609FC, 32'hFEEAF50F, 32'hFE07ED03, 32'hFF17FE0D, 
    /* (5, 0) */	    32'hE51509FC, 32'hFEEBF50E, 32'hFE06EE03, 32'hFF16FE0C, 
    /* (6, 0) */	    32'hE61409FC, 32'hFEEBF60E, 32'hFE06EE03, 32'hFF15FE0C, 
    /* (7, 0) */	    32'hE71408FC, 32'hFEECF60D, 32'hFE06EF02, 32'hFF14FE0B, 
    /* (8, 0) */	    32'hE81308FD, 32'hFEEDF70D, 32'hFE06F002, 32'hFF13FE0B, 
    /* (9, 0) */	    32'hE91208FD, 32'hFEEEF70C, 32'hFE05F002, 32'hFF13FE0A, 
    /* (10, 0) */	    32'hEA1107FD, 32'hFEEFF70C, 32'hFE05F102, 32'hFF12FE0A, 
    /* (11, 0) */	    32'hEB1107FD, 32'hFEEFF80B, 32'hFE05F202, 32'hFF11FE09, 
    /* (12, 0) */	    32'hEC1007FD, 32'hFEF0F80B, 32'hFE05F202, 32'hFF10FE09, 
    /* (13, 0) */	    32'hED0F06FD, 32'hFFF1F90A, 32'hFE04F302, 32'hFF0FFE09, 
    /* (14, 0) */	    32'hEE0E06FD, 32'hFFF2F90A, 32'hFE04F402, 32'hFF0FFF08, 
    /* (15, 0) */	    32'hEF0D06FE, 32'hFFF3F909, 32'hFF04F402, 32'hFF0EFF08, 
    /* (16, 0) */	    32'hF00D05FE, 32'hFFF3FA08, 32'hFF04F502, 32'hFF0DFF07, 
    /* (17, 0) */	    32'hF10C05FE, 32'hFFF4FA08, 32'hFF04F601, 32'hFF0CFF07, 
    /* (18, 0) */	    32'hF20B05FE, 32'hFFF5FA07, 32'hFF03F601, 32'hFF0BFF06, 
    /* (19, 0) */	    32'hF30A04FE, 32'hFFF6FB07, 32'hFF03F701, 32'hFF0BFF06, 
    /* (20, 0) */	    32'hF40904FE, 32'hFFF6FB06, 32'hFF03F801, 32'hFF0AFF05, 
    /* (21, 0) */	    32'hF50904FE, 32'hFFF7FC06, 32'hFF03F901, 32'hFF09FF05, 
    /* (22, 0) */	    32'hF60803FF, 32'hFFF8FC05, 32'hFF02F901, 32'hFF08FF05, 
    /* (23, 0) */	    32'hF70703FF, 32'hFFF9FC05, 32'hFF02FA01, 32'h0007FF04, 
    /* (24, 0) */	    32'hF80603FF, 32'hFFFAFD04, 32'hFF02FB01, 32'h0006FF04, 
    /* (25, 0) */	    32'hF90602FF, 32'hFFFAFD04, 32'hFF02FB01, 32'h0006FF03, 
    /* (26, 0) */	    32'hFA0502FF, 32'h00FBFE03, 32'hFF01FC01, 32'h00050003, 
    /* (27, 0) */	    32'hFB0402FF, 32'h00FCFE03, 32'h0001FD00, 32'h00040002, 
    /* (28, 0) */	    32'hFC0301FF, 32'h00FDFE02, 32'h0001FD00, 32'h00030002, 
    /* (29, 0) */	    32'hFD020100, 32'h00FEFF02, 32'h0001FE00, 32'h00020001, 
    /* (30, 0) */	    32'hFE020100, 32'h00FEFF01, 32'h0000FF00, 32'h00020001, 
    /* (31, 0) */	    32'hFF010000, 32'h00FF0001, 32'h0000FF00, 32'h00010000, 
    /* (32, 0) */	    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
    /* (33, 0) */	    32'h01FF0000, 32'h000100FF, 32'h00000100, 32'h00FF0000, 
    /* (34, 0) */	    32'h02FEFF00, 32'h000201FF, 32'h00000100, 32'h00FE00FF, 
    /* (35, 0) */	    32'h03FEFF00, 32'h000201FE, 32'h00FF0200, 32'h00FE00FF, 
    /* (36, 0) */	    32'h04FDFF01, 32'h000302FE, 32'h00FF0300, 32'h00FD00FE, 
    /* (37, 0) */	    32'h05FCFE01, 32'h000402FD, 32'h00FF0300, 32'h00FC00FE, 
    /* (38, 0) */	    32'h06FBFE01, 32'h000502FD, 32'h01FF04FF, 32'h00FB00FD, 
    /* (39, 0) */	    32'h07FAFE01, 32'h010603FC, 32'h01FE05FF, 32'h00FA01FD, 
    /* (40, 0) */	    32'h08FAFD01, 32'h010603FC, 32'h01FE05FF, 32'h00FA01FC, 
    /* (41, 0) */	    32'h09F9FD01, 32'h010704FB, 32'h01FE06FF, 32'h00F901FC, 
    /* (42, 0) */	    32'h0AF8FD01, 32'h010804FB, 32'h01FE07FF, 32'h01F801FB, 
    /* (43, 0) */	    32'h0BF7FC02, 32'h010904FA, 32'h01FD07FF, 32'h01F701FB, 
    /* (44, 0) */	    32'h0CF7FC02, 32'h010A05FA, 32'h01FD08FF, 32'h01F601FB, 
    /* (45, 0) */	    32'h0DF6FC02, 32'h010A05F9, 32'h01FD09FF, 32'h01F501FA, 
    /* (46, 0) */	    32'h0EF5FB02, 32'h010B06F9, 32'h01FD0AFF, 32'h01F501FA, 
    /* (47, 0) */	    32'h0FF4FB02, 32'h010C06F8, 32'h01FC0AFF, 32'h01F401F9, 
    /* (48, 0) */	    32'h10F3FB02, 32'h010D06F8, 32'h01FC0BFE, 32'h01F301F9, 
    /* (49, 0) */	    32'h11F3FA02, 32'h010D07F7, 32'h01FC0CFE, 32'h01F201F8, 
    /* (50, 0) */	    32'h12F2FA03, 32'h010E07F6, 32'h02FC0CFE, 32'h01F101F8, 
    /* (51, 0) */	    32'h13F1FA03, 32'h010F07F6, 32'h02FC0DFE, 32'h01F102F7, 
    /* (52, 0) */	    32'h14F0F903, 32'h021008F5, 32'h02FB0EFE, 32'h01F002F7, 
    /* (53, 0) */	    32'h15EFF903, 32'h021108F5, 32'h02FB0EFE, 32'h01EF02F7, 
    /* (54, 0) */	    32'h16EFF903, 32'h021109F4, 32'h02FB0FFE, 32'h01EE02F6, 
    /* (55, 0) */	    32'h17EEF803, 32'h021209F4, 32'h02FB10FE, 32'h01ED02F6, 
    /* (56, 0) */	    32'h18EDF803, 32'h021309F3, 32'h02FA10FE, 32'h01ED02F5, 
    /* (57, 0) */	    32'h19ECF804, 32'h02140AF3, 32'h02FA11FE, 32'h01EC02F5, 
    /* (58, 0) */	    32'h1AECF704, 32'h02150AF2, 32'h02FA12FD, 32'h01EB02F4, 
    /* (59, 0) */	    32'h1BEBF704, 32'h02150BF2, 32'h02FA12FD, 32'h01EA02F4, 
    /* (60, 0) */	    32'h1BEAF704, 32'h02160BF1, 32'h02F913FD, 32'h01E902F3, 
    /* (61, 0) */	    32'h1CE9F604, 32'h02170BF1, 32'h02F914FD, 32'h01E902F3, 
    /* (62, 0) */	    32'h1DE8F604, 32'h02180CF0, 32'h03F914FD, 32'h02E802F2, 
    /* (63, 0) */	    32'h1EE8F504, 32'h02190CF0, 32'h03F915FD, 32'h02E703F2, 
    /* (64, 0) */	    32'h12DFF409, 32'hE9ED43F5, 32'h50FF08F8, 32'h32D0F3F2, 
    /* (65, 0) */	    32'h12E1F409, 32'hEAED41F5, 32'h4DFF08F8, 32'h30D1F4F2, 
    /* (66, 0) */	    32'h11E2F509, 32'hEBEE3FF5, 32'h4BFF07F8, 32'h2ED3F4F3, 
    /* (67, 0) */	    32'h11E3F508, 32'hEBEE3DF6, 32'h48FF07F8, 32'h2DD4F4F3, 
    /* (68, 0) */	    32'h10E4F608, 32'hECEF3BF6, 32'h46FF07F9, 32'h2BD6F5F4, 
    /* (69, 0) */	    32'h0FE5F608, 32'hEDF039F6, 32'h43FF07F9, 32'h2AD7F5F4, 
    /* (70, 0) */	    32'h0FE6F607, 32'hEDF036F7, 32'h41FF06F9, 32'h28D9F6F5, 
    /* (71, 0) */	    32'h0EE7F707, 32'hEEF134F7, 32'h3EFF06F9, 32'h27DAF6F5, 
    /* (72, 0) */	    32'h0EE8F707, 32'hEFF132F7, 32'h3CFF06FA, 32'h25DCF6F6, 
    /* (73, 0) */	    32'h0DE9F707, 32'hF0F230F8, 32'h39FF06FA, 32'h24DDF7F6, 
    /* (74, 0) */	    32'h0DEAF806, 32'hF0F32EF8, 32'h37FF05FA, 32'h22DFF7F6, 
    /* (75, 0) */	    32'h0CEBF806, 32'hF1F32CF8, 32'h340005FA, 32'h21E0F8F7, 
    /* (76, 0) */	    32'h0BECF906, 32'hF2F42AF9, 32'h320005FB, 32'h1FE2F8F7, 
    /* (77, 0) */	    32'h0BEDF905, 32'hF2F428F9, 32'h2F0005FB, 32'h1DE3F8F8, 
    /* (78, 0) */	    32'h0AEEF905, 32'hF3F526FA, 32'h2D0004FB, 32'h1CE5F9F8, 
    /* (79, 0) */	    32'h0AEFFA05, 32'hF4F624FA, 32'h2A0004FB, 32'h1AE6F9F9, 
    /* (80, 0) */	    32'h09F0FA05, 32'hF5F622FA, 32'h280004FC, 32'h19E8FAF9, 
    /* (81, 0) */	    32'h09F1FA04, 32'hF5F71FFB, 32'h250004FC, 32'h17E9FAF9, 
    /* (82, 0) */	    32'h08F2FB04, 32'hF6F71DFB, 32'h230003FC, 32'h16EBFAFA, 
    /* (83, 0) */	    32'h07F3FB04, 32'hF7F81BFB, 32'h200003FD, 32'h14ECFBFA, 
    /* (84, 0) */	    32'h07F4FC03, 32'hF7F919FC, 32'h1E0003FD, 32'h13EEFBFB, 
    /* (85, 0) */	    32'h06F5FC03, 32'hF8F917FC, 32'h1B0003FD, 32'h11EFFCFB, 
    /* (86, 0) */	    32'h06F6FC03, 32'hF9FA15FC, 32'h190002FD, 32'h0FF1FCFC, 
    /* (87, 0) */	    32'h05F7FD03, 32'hFAFB13FD, 32'h160002FE, 32'h0EF2FCFC, 
    /* (88, 0) */	    32'h05F8FD02, 32'hFAFB11FD, 32'h140002FE, 32'h0CF4FDFD, 
    /* (89, 0) */	    32'h04F9FD02, 32'hFBFC0FFD, 32'h110002FE, 32'h0BF5FDFD, 
    /* (90, 0) */	    32'h03FAFE02, 32'hFCFC0DFE, 32'h0F0001FE, 32'h09F7FEFD, 
    /* (91, 0) */	    32'h03FBFE01, 32'hFCFD0AFE, 32'h0C0001FF, 32'h08F8FEFE, 
    /* (92, 0) */	    32'h02FCFF01, 32'hFDFE08FF, 32'h0A0001FF, 32'h06FAFEFE, 
    /* (93, 0) */	    32'h02FDFF01, 32'hFEFE06FF, 32'h070001FF, 32'h05FBFFFF, 
    /* (94, 0) */	    32'h01FEFF01, 32'hFFFF04FF, 32'h050000FF, 32'h03FDFFFF, 
    /* (95, 0) */	    32'h01FF0000, 32'hFFFF0200, 32'h02000000, 32'h02FE0000, 
    /* (96, 0) */	    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
    /* (97, 0) */	    32'hFF010000, 32'h0101FE00, 32'hFE000000, 32'hFE020000, 
    /* (98, 0) */	    32'hFF0201FF, 32'h0101FC01, 32'hFB000001, 32'hFD030101, 
    /* (99, 0) */	    32'hFE0301FF, 32'h0202FA01, 32'hF900FF01, 32'hFB050101, 
    /* (100, 0) */	    32'hFE0401FF, 32'h0302F801, 32'hF600FF01, 32'hFA060202, 
    /* (101, 0) */	    32'hFD0502FF, 32'h0403F602, 32'hF400FF01, 32'hF8080202, 
    /* (102, 0) */	    32'hFD0602FE, 32'h0404F302, 32'hF100FF02, 32'hF7090203, 
    /* (103, 0) */	    32'hFC0703FE, 32'h0504F103, 32'hEF00FE02, 32'hF50B0303, 
    /* (104, 0) */	    32'hFB0803FE, 32'h0605EF03, 32'hEC00FE02, 32'hF40C0303, 
    /* (105, 0) */	    32'hFB0903FD, 32'h0605ED03, 32'hEA00FE02, 32'hF20E0404, 
    /* (106, 0) */	    32'hFA0A04FD, 32'h0706EB04, 32'hE700FE03, 32'hF10F0404, 
    /* (107, 0) */	    32'hFA0B04FD, 32'h0807E904, 32'hE500FD03, 32'hEF110405, 
    /* (108, 0) */	    32'hF90C04FD, 32'h0907E704, 32'hE200FD03, 32'hED120505, 
    /* (109, 0) */	    32'hF90D05FC, 32'h0908E505, 32'hE000FD03, 32'hEC140506, 
    /* (110, 0) */	    32'hF80E05FC, 32'h0A09E305, 32'hDD00FD04, 32'hEA150606, 
    /* (111, 0) */	    32'hF70F06FC, 32'h0B09E105, 32'hDB00FC04, 32'hE9170607, 
    /* (112, 0) */	    32'hF71006FB, 32'h0B0ADE06, 32'hD800FC04, 32'hE7180607, 
    /* (113, 0) */	    32'hF61106FB, 32'h0C0ADC06, 32'hD600FC05, 32'hE61A0707, 
    /* (114, 0) */	    32'hF61207FB, 32'h0D0BDA06, 32'hD300FC05, 32'hE41B0708, 
    /* (115, 0) */	    32'hF51307FB, 32'h0E0CD807, 32'hD100FB05, 32'hE31D0808, 
    /* (116, 0) */	    32'hF51407FA, 32'h0E0CD607, 32'hCE00FB05, 32'hE11E0809, 
    /* (117, 0) */	    32'hF41508FA, 32'h0F0DD408, 32'hCC00FB06, 32'hDF200809, 
    /* (118, 0) */	    32'hF31608FA, 32'h100DD208, 32'hC901FB06, 32'hDE21090A, 
    /* (119, 0) */	    32'hF31709F9, 32'h100ED008, 32'hC701FA06, 32'hDC23090A, 
    /* (120, 0) */	    32'hF21809F9, 32'h110FCE09, 32'hC401FA06, 32'hDB240A0A, 
    /* (121, 0) */	    32'hF21909F9, 32'h120FCC09, 32'hC201FA07, 32'hD9260A0B, 
    /* (122, 0) */	    32'hF11A0AF9, 32'h1310CA09, 32'hBF01FA07, 32'hD8270A0B, 
    /* (123, 0) */	    32'hF11B0AF8, 32'h1310C70A, 32'hBD01F907, 32'hD6290B0C, 
    /* (124, 0) */	    32'hF01C0AF8, 32'h1411C50A, 32'hBA01F907, 32'hD52A0B0C, 
    /* (125, 0) */	    32'hEF1D0BF8, 32'h1512C30A, 32'hB801F908, 32'hD32C0C0D, 
    /* (126, 0) */	    32'hEF1E0BF7, 32'h1512C10B, 32'hB501F908, 32'hD22D0C0D, 
    /* (127, 0) */	    32'hEE1F0CF7, 32'h1613BF0B, 32'hB301F808, 32'hD02F0C0E, 
    /* (128, 0) */	    32'h37FB39FA, 32'h38807FF6, 32'hD6F0E4ED, 32'hE2DA12C9, 
    /* (129, 0) */	    32'h36FB37FA, 32'h36847BF6, 32'hD7F0E5EE, 32'hE3DB11CB, 
    /* (130, 0) */	    32'h34FB35FA, 32'h348878F6, 32'hD9F1E6EE, 32'hE4DC11CD, 
    /* (131, 0) */	    32'h32FB33FA, 32'h328C74F7, 32'hDAF1E7EF, 32'hE5DE10CE, 
    /* (132, 0) */	    32'h30FB32FB, 32'h319070F7, 32'hDBF2E8EF, 32'hE6DF10D0, 
    /* (133, 0) */	    32'h2FFC30FB, 32'h2F946CF7, 32'hDDF2E9F0, 32'hE7E00FD2, 
    /* (134, 0) */	    32'h2DFC2EFB, 32'h2D9868F8, 32'hDEF3EAF1, 32'hE8E10ED3, 
    /* (135, 0) */	    32'h2BFC2CFB, 32'h2B9C64F8, 32'hDFF3EAF1, 32'hE9E20ED5, 
    /* (136, 0) */	    32'h29FC2BFB, 32'h2AA060F8, 32'hE1F4EBF2, 32'hEAE40DD7, 
    /* (137, 0) */	    32'h28FC29FC, 32'h28A45CF9, 32'hE2F4ECF2, 32'hEBE50DD9, 
    /* (138, 0) */	    32'h26FC27FC, 32'h26A858F9, 32'hE3F5EDF3, 32'hECE60CDA, 
    /* (139, 0) */	    32'h24FD25FC, 32'h24AC54F9, 32'hE5F5EEF4, 32'hEDE70CDC, 
    /* (140, 0) */	    32'h23FD23FC, 32'h23B050FA, 32'hE6F6EFF4, 32'hEEE80BDE, 
    /* (141, 0) */	    32'h21FD22FC, 32'h21B44CFA, 32'hE7F6F0F5, 32'hEEEA0BDF, 
    /* (142, 0) */	    32'h1FFD20FD, 32'h1FB848FA, 32'hE8F7F0F5, 32'hEFEB0AE1, 
    /* (143, 0) */	    32'h1DFD1EFD, 32'h1EBC44FB, 32'hEAF7F1F6, 32'hF0EC09E3, 
    /* (144, 0) */	    32'h1CFD1CFD, 32'h1CC040FB, 32'hEBF8F2F7, 32'hF1ED09E5, 
    /* (145, 0) */	    32'h1AFE1BFD, 32'h1AC43CFB, 32'hECF8F3F7, 32'hF2EE08E6, 
    /* (146, 0) */	    32'h18FE19FD, 32'h18C838FB, 32'hEEF9F4F8, 32'hF3EF08E8, 
    /* (147, 0) */	    32'h16FE17FD, 32'h17CC34FC, 32'hEFF9F5F8, 32'hF4F107EA, 
    /* (148, 0) */	    32'h15FE15FE, 32'h15D030FC, 32'hF0FAF6F9, 32'hF5F207EB, 
    /* (149, 0) */	    32'h13FE13FE, 32'h13D42CFC, 32'hF2FAF7F9, 32'hF6F306ED, 
    /* (150, 0) */	    32'h11FE12FE, 32'h11D828FD, 32'hF3FBF7FA, 32'hF7F406EF, 
    /* (151, 0) */	    32'h10FF10FE, 32'h10DC24FD, 32'hF4FBF8FB, 32'hF8F505F1, 
    /* (152, 0) */	    32'h0EFF0EFE, 32'h0EE020FD, 32'hF6FCF9FB, 32'hF9F704F2, 
    /* (153, 0) */	    32'h0CFF0CFF, 32'h0CE41CFE, 32'hF7FCFAFC, 32'hFAF804F4, 
    /* (154, 0) */	    32'h0AFF0BFF, 32'h0AE818FE, 32'hF8FDFBFC, 32'hFAF903F6, 
    /* (155, 0) */	    32'h09FF09FF, 32'h09EC14FE, 32'hF9FDFCFD, 32'hFBFA03F7, 
    /* (156, 0) */	    32'h07FF07FF, 32'h07F010FF, 32'hFBFEFDFE, 32'hFCFB02F9, 
    /* (157, 0) */	    32'h050005FF, 32'h05F40CFF, 32'hFCFEFDFE, 32'hFDFC02FB, 
    /* (158, 0) */	    32'h03000400, 32'h03F808FF, 32'hFDFFFEFF, 32'hFEFE01FD, 
    /* (159, 0) */	    32'h02000200, 32'h02FC0400, 32'hFFFFFFFF, 32'hFFFF01FE, 
    /* (160, 0) */	    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
    /* (161, 0) */	    32'hFE00FE00, 32'hFE04FC00, 32'h01010101, 32'h0101FF02, 
    /* (162, 0) */	    32'hFD00FC00, 32'hFD08F801, 32'h03010201, 32'h0202FF03, 
    /* (163, 0) */	    32'hFB00FB01, 32'hFB0CF401, 32'h04020302, 32'h0304FE05, 
    /* (164, 0) */	    32'hF901F901, 32'hF910F001, 32'h05020302, 32'h0405FE07, 
    /* (165, 0) */	    32'hF701F701, 32'hF714EC02, 32'h07030403, 32'h0506FD09, 
    /* (166, 0) */	    32'hF601F501, 32'hF618E802, 32'h08030504, 32'h0607FD0A, 
    /* (167, 0) */	    32'hF401F401, 32'hF41CE402, 32'h09040604, 32'h0608FC0C, 
    /* (168, 0) */	    32'hF201F202, 32'hF220E003, 32'h0A040705, 32'h0709FC0E, 
    /* (169, 0) */	    32'hF001F002, 32'hF024DC03, 32'h0C050805, 32'h080BFB0F, 
    /* (170, 0) */	    32'hEF02EE02, 32'hEF28D803, 32'h0D050906, 32'h090CFA11, 
    /* (171, 0) */	    32'hED02ED02, 32'hED2CD404, 32'h0E060907, 32'h0A0DFA13, 
    /* (172, 0) */	    32'hEB02EB02, 32'hEB30D004, 32'h10060A07, 32'h0B0EF915, 
    /* (173, 0) */	    32'hEA02E903, 32'hE934CC04, 32'h11070B08, 32'h0C0FF916, 
    /* (174, 0) */	    32'hE802E703, 32'hE838C805, 32'h12070C08, 32'h0D11F818, 
    /* (175, 0) */	    32'hE602E503, 32'hE63CC405, 32'h14080D09, 32'h0E12F81A, 
    /* (176, 0) */	    32'hE403E403, 32'hE440C005, 32'h15080E09, 32'h0F13F71B, 
    /* (177, 0) */	    32'hE303E203, 32'hE244BC05, 32'h16090F0A, 32'h1014F71D, 
    /* (178, 0) */	    32'hE103E003, 32'hE148B806, 32'h1809100B, 32'h1115F61F, 
    /* (179, 0) */	    32'hDF03DE04, 32'hDF4CB406, 32'h190A100B, 32'h1216F521, 
    /* (180, 0) */	    32'hDD03DD04, 32'hDD50B006, 32'h1A0A110C, 32'h1218F522, 
    /* (181, 0) */	    32'hDC03DB04, 32'hDC54AC07, 32'h1B0B120C, 32'h1319F424, 
    /* (182, 0) */	    32'hDA04D904, 32'hDA58A807, 32'h1D0B130D, 32'h141AF426, 
    /* (183, 0) */	    32'hD804D704, 32'hD85CA407, 32'h1E0C140E, 32'h151BF327, 
    /* (184, 0) */	    32'hD704D505, 32'hD660A008, 32'h1F0C150E, 32'h161CF329, 
    /* (185, 0) */	    32'hD504D405, 32'hD5649C08, 32'h210D160F, 32'h171EF22B, 
    /* (186, 0) */	    32'hD304D205, 32'hD3689808, 32'h220D160F, 32'h181FF22D, 
    /* (187, 0) */	    32'hD104D005, 32'hD16C9409, 32'h230E1710, 32'h1920F12E, 
    /* (188, 0) */	    32'hD005CE05, 32'hCF709009, 32'h250E1811, 32'h1A21F030, 
    /* (189, 0) */	    32'hCE05CD06, 32'hCE748C09, 32'h260F1911, 32'h1B22F032, 
    /* (190, 0) */	    32'hCC05CB06, 32'hCC78880A, 32'h270F1A12, 32'h1C24EF33, 
    /* (191, 0) */	    32'hCA05C906, 32'hCA7C850A, 32'h29101B12, 32'h1D25EF35, 
    /* (192, 0) */	    32'hE8F7FB2E, 32'h180C10F4, 32'h15FA23F6, 32'hFCD2FFFF, 
    /* (193, 0) */	    32'hE8F7FB2C, 32'h180C0FF5, 32'h14FB22F6, 32'hFCD3FFFF, 
    /* (194, 0) */	    32'hE9F8FB2B, 32'h170B0FF5, 32'h14FB21F6, 32'hFDD5FFFF, 
    /* (195, 0) */	    32'hEAF8FB2A, 32'h160B0EF5, 32'h13FB20F7, 32'hFDD6FF00, 
    /* (196, 0) */	    32'hEBF8FB28, 32'h150B0EF6, 32'h12FB1FF7, 32'hFDD8FF00, 
    /* (197, 0) */	    32'hEBF8FC27, 32'h140A0DF6, 32'h12FB1EF7, 32'hFDD9FF00, 
    /* (198, 0) */	    32'hECF9FC25, 32'h140A0DF6, 32'h11FB1DF8, 32'hFDDAFF00, 
    /* (199, 0) */	    32'hEDF9FC24, 32'h13090CF7, 32'h10FC1CF8, 32'hFDDCFF00, 
    /* (200, 0) */	    32'hEEF9FC22, 32'h12090CF7, 32'h10FC1BF8, 32'hFDDDFF00, 
    /* (201, 0) */	    32'hEFFAFC21, 32'h11090BF8, 32'h0FFC19F9, 32'hFDDFFF00, 
    /* (202, 0) */	    32'hEFFAFC1F, 32'h11080BF8, 32'h0EFC18F9, 32'hFDE0FF00, 
    /* (203, 0) */	    32'hF0FAFD1E, 32'h10080AF8, 32'h0EFC17F9, 32'hFEE2FF00, 
    /* (204, 0) */	    32'hF1FAFD1D, 32'h0F080AF9, 32'h0DFD16FA, 32'hFEE3FF00, 
    /* (205, 0) */	    32'hF2FBFD1B, 32'h0E0709F9, 32'h0CFD15FA, 32'hFEE5FF00, 
    /* (206, 0) */	    32'hF2FBFD1A, 32'h0E0709F9, 32'h0CFD14FA, 32'hFEE6FF00, 
    /* (207, 0) */	    32'hF3FBFD18, 32'h0D0608FA, 32'h0BFD13FB, 32'hFEE7FF00, 
    /* (208, 0) */	    32'hF4FBFD17, 32'h0C0608FA, 32'h0AFD12FB, 32'hFEE9FF00, 
    /* (209, 0) */	    32'hF5FCFE15, 32'h0B0607FA, 32'h0AFD11FB, 32'hFEEAFF00, 
    /* (210, 0) */	    32'hF5FCFE14, 32'h0B0507FB, 32'h09FE0FFC, 32'hFEECFF00, 
    /* (211, 0) */	    32'hF6FCFE13, 32'h0A0506FB, 32'h08FE0EFC, 32'hFEED0000, 
    /* (212, 0) */	    32'hF7FDFE11, 32'h090506FC, 32'h08FE0DFC, 32'hFFEF0000, 
    /* (213, 0) */	    32'hF8FDFE10, 32'h080405FC, 32'h07FE0CFC, 32'hFFF00000, 
    /* (214, 0) */	    32'hF8FDFE0E, 32'h080405FC, 32'h07FE0BFD, 32'hFFF20000, 
    /* (215, 0) */	    32'hF9FDFF0D, 32'h070304FD, 32'h06FE0AFD, 32'hFFF30000, 
    /* (216, 0) */	    32'hFAFEFF0B, 32'h060304FD, 32'h05FF09FD, 32'hFFF40000, 
    /* (217, 0) */	    32'hFBFEFF0A, 32'h050303FD, 32'h05FF08FE, 32'hFFF60000, 
    /* (218, 0) */	    32'hFBFEFF09, 32'h050203FE, 32'h04FF07FE, 32'hFFF70000, 
    /* (219, 0) */	    32'hFCFFFF07, 32'h040202FE, 32'h03FF06FE, 32'hFFF90000, 
    /* (220, 0) */	    32'hFDFFFF06, 32'h030202FF, 32'h03FF04FF, 32'h00FA0000, 
    /* (221, 0) */	    32'hFEFF0004, 32'h020101FF, 32'h02FF03FF, 32'h00FC0000, 
    /* (222, 0) */	    32'hFEFF0003, 32'h020101FF, 32'h010002FF, 32'h00FD0000, 
    /* (223, 0) */	    32'hFF000001, 32'h01000000, 32'h01000100, 32'h00FF0000, 
    /* (224, 0) */	    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
    /* (225, 0) */	    32'h010000FF, 32'hFF000000, 32'hFF00FF00, 32'h00010000, 
    /* (226, 0) */	    32'h020100FD, 32'hFEFFFF01, 32'hFF00FE01, 32'h00030000, 
    /* (227, 0) */	    32'h020100FC, 32'hFEFFFF01, 32'hFE01FD01, 32'h00040000, 
    /* (228, 0) */	    32'h030101FA, 32'hFDFEFE01, 32'hFD01FC01, 32'h00060000, 
    /* (229, 0) */	    32'h040101F9, 32'hFCFEFE02, 32'hFD01FA02, 32'h01070000, 
    /* (230, 0) */	    32'h050201F7, 32'hFBFEFD02, 32'hFC01F902, 32'h01090000, 
    /* (231, 0) */	    32'h050201F6, 32'hFBFDFD03, 32'hFB01F802, 32'h010A0000, 
    /* (232, 0) */	    32'h060201F5, 32'hFAFDFC03, 32'hFB01F703, 32'h010C0000, 
    /* (233, 0) */	    32'h070301F3, 32'hF9FDFC03, 32'hFA02F603, 32'h010D0000, 
    /* (234, 0) */	    32'h080302F2, 32'hF8FCFB04, 32'hF902F503, 32'h010E0000, 
    /* (235, 0) */	    32'h080302F0, 32'hF8FCFB04, 32'hF902F404, 32'h01100000, 
    /* (236, 0) */	    32'h090302EF, 32'hF7FBFA04, 32'hF802F304, 32'h01110000, 
    /* (237, 0) */	    32'h0A0402ED, 32'hF6FBFA05, 32'hF802F204, 32'h02130000, 
    /* (238, 0) */	    32'h0B0402EC, 32'hF5FBF905, 32'hF702F104, 32'h02140100, 
    /* (239, 0) */	    32'h0B0402EB, 32'hF5FAF906, 32'hF603EF05, 32'h02160100, 
    /* (240, 0) */	    32'h0C0503E9, 32'hF4FAF806, 32'hF603EE05, 32'h02170100, 
    /* (241, 0) */	    32'h0D0503E8, 32'hF3FAF806, 32'hF503ED05, 32'h02190100, 
    /* (242, 0) */	    32'h0E0503E6, 32'hF2F9F707, 32'hF403EC06, 32'h021A0100, 
    /* (243, 0) */	    32'h0E0503E5, 32'hF2F9F707, 32'hF403EB06, 32'h021B0100, 
    /* (244, 0) */	    32'h0F0603E3, 32'hF1F8F607, 32'hF303EA06, 32'h021D0100, 
    /* (245, 0) */	    32'h100603E2, 32'hF0F8F608, 32'hF204E907, 32'h021E0100, 
    /* (246, 0) */	    32'h110604E1, 32'hEFF8F508, 32'hF204E807, 32'h03200100, 
    /* (247, 0) */	    32'h110604DF, 32'hEFF7F508, 32'hF104E707, 32'h03210100, 
    /* (248, 0) */	    32'h120704DE, 32'hEEF7F409, 32'hF004E508, 32'h03230100, 
    /* (249, 0) */	    32'h130704DC, 32'hEDF7F409, 32'hF004E408, 32'h03240100, 
    /* (250, 0) */	    32'h140704DB, 32'hECF6F30A, 32'hEF05E308, 32'h03260100, 
    /* (251, 0) */	    32'h150804D9, 32'hECF6F30A, 32'hEE05E209, 32'h03270100, 
    /* (252, 0) */	    32'h150805D8, 32'hEBF5F20A, 32'hEE05E109, 32'h03280100, 
    /* (253, 0) */	    32'h160805D6, 32'hEAF5F20B, 32'hED05E009, 32'h032A0100, 
    /* (254, 0) */	    32'h170805D5, 32'hE9F5F10B, 32'hEC05DF0A, 32'h032B0101, 
    /* (255, 0) */	    32'h180905D4, 32'hE8F4F10B, 32'hEC05DE0A, 32'h042D0101, 
    /* (256, 0) */	    32'h7F7FCFCF, 32'hFEDEA3B7, 32'h9F01D1B2, 32'hCF07337F, 
    /* (257, 0) */	    32'h7F7BD1D1, 32'hFEDFA6B9, 32'hA201D3B4, 32'hD006317C, 
    /* (258, 0) */	    32'h7F77D2D2, 32'hFFE0A9BB, 32'hA501D4B7, 32'hD2063078, 
    /* (259, 0) */	    32'h7C74D4D4, 32'hFFE1ACBE, 32'hA801D6B9, 32'hD3062E74, 
    /* (260, 0) */	    32'h7870D5D5, 32'hFFE2AEC0, 32'hAB01D7BC, 32'hD5062D70, 
    /* (261, 0) */	    32'h746CD7D7, 32'hFFE3B1C2, 32'hAE01D9BE, 32'hD6062B6C, 
    /* (262, 0) */	    32'h6F68D8D8, 32'hFFE4B4C5, 32'hB101DAC1, 32'hD8052968, 
    /* (263, 0) */	    32'h6B64DADA, 32'hFFE5B7C7, 32'hB401DCC3, 32'hD9052864, 
    /* (264, 0) */	    32'h6760DBDB, 32'hFFE6BAC9, 32'hB701DDC6, 32'hDB052660, 
    /* (265, 0) */	    32'h635CDDDD, 32'hFFE8BDCB, 32'hBA01DEC8, 32'hDD05255C, 
    /* (266, 0) */	    32'h5E58DEDE, 32'hFFE9C0CE, 32'hBD01E0CA, 32'hDE052358, 
    /* (267, 0) */	    32'h5A54E0E0, 32'hFFEAC3D0, 32'hC101E1CD, 32'hE0042154, 
    /* (268, 0) */	    32'h5650E1E1, 32'hFFEBC6D2, 32'hC401E3CF, 32'hE1042050, 
    /* (269, 0) */	    32'h514CE3E3, 32'hFFECC9D5, 32'hC701E4D2, 32'hE3041E4C, 
    /* (270, 0) */	    32'h4D48E5E5, 32'hFFEDCCD7, 32'hCA01E6D4, 32'hE4041D48, 
    /* (271, 0) */	    32'h4944E6E6, 32'hFFEECED9, 32'hCD01E7D7, 32'hE6041B44, 
    /* (272, 0) */	    32'h4540E8E8, 32'hFFEFD1DB, 32'hD001E9D9, 32'hE7031940, 
    /* (273, 0) */	    32'h403CE9E9, 32'hFFF0D4DE, 32'hD301EADB, 32'hE903183C, 
    /* (274, 0) */	    32'h3C38EBEB, 32'hFFF1D7E0, 32'hD601ECDE, 32'hEA031638, 
    /* (275, 0) */	    32'h3834ECEC, 32'hFFF2DAE2, 32'hD901EDE0, 32'hEC031534, 
    /* (276, 0) */	    32'h3330EEEE, 32'hFFF3DDE5, 32'hDC01EEE3, 32'hEE021330, 
    /* (277, 0) */	    32'h2F2CEFEF, 32'hFFF4E0E7, 32'hDF01F0E5, 32'hEF02122C, 
    /* (278, 0) */	    32'h2B28F1F1, 32'h00F5E3E9, 32'hE200F1E8, 32'hF1021028, 
    /* (279, 0) */	    32'h2724F2F2, 32'h00F6E6EB, 32'hE500F3EA, 32'hF2020E24, 
    /* (280, 0) */	    32'h2220F4F4, 32'h00F7E9EE, 32'hE800F4ED, 32'hF4020D20, 
    /* (281, 0) */	    32'h1E1CF5F5, 32'h00F9ECF0, 32'hEB00F6EF, 32'hF5010B1C, 
    /* (282, 0) */	    32'h1A18F7F7, 32'h00FAEFF2, 32'hEE00F7F1, 32'hF7010A18, 
    /* (283, 0) */	    32'h1514F8F8, 32'h00FBF1F5, 32'hF100F9F4, 32'hF8010814, 
    /* (284, 0) */	    32'h1110FAFA, 32'h00FCF4F7, 32'hF400FAF6, 32'hFA010610, 
    /* (285, 0) */	    32'h0D0CFBFB, 32'h00FDF7F9, 32'hF700FCF9, 32'hFB01050C, 
    /* (286, 0) */	    32'h0908FDFD, 32'h00FEFAFB, 32'hFA00FDFB, 32'hFD000308, 
    /* (287, 0) */	    32'h0404FEFE, 32'h00FFFDFE, 32'hFD00FFFE, 32'hFE000204, 
    /* (288, 0) */	    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
    /* (289, 0) */	    32'hFCFC0202, 32'h00010302, 32'h03000102, 32'h0200FEFC, 
    /* (290, 0) */	    32'hF7F80303, 32'h00020605, 32'h06000305, 32'h0300FDF8, 
    /* (291, 0) */	    32'hF3F40505, 32'h00030907, 32'h09000407, 32'h05FFFBF4, 
    /* (292, 0) */	    32'hEFF00606, 32'h00040C09, 32'h0C00060A, 32'h06FFFAF0, 
    /* (293, 0) */	    32'hEBEC0808, 32'h00050F0B, 32'h0F00070C, 32'h08FFF8EC, 
    /* (294, 0) */	    32'hE6E80909, 32'h0006110E, 32'h1200090F, 32'h09FFF6E8, 
    /* (295, 0) */	    32'hE2E40B0B, 32'h00071410, 32'h15000A11, 32'h0BFFF5E4, 
    /* (296, 0) */	    32'hDEE00C0C, 32'h00091712, 32'h18000C13, 32'h0CFEF3E0, 
    /* (297, 0) */	    32'hD9DC0E0E, 32'h000A1A15, 32'h1B000D16, 32'h0EFEF2DC, 
    /* (298, 0) */	    32'hD5D80F0F, 32'h000B1D17, 32'h1E000F18, 32'h0FFEF0D8, 
    /* (299, 0) */	    32'hD1D41111, 32'h010C2019, 32'h21FF101B, 32'h11FEEED4, 
    /* (300, 0) */	    32'hCDD01212, 32'h010D231B, 32'h24FF121D, 32'h12FEEDD0, 
    /* (301, 0) */	    32'hC8CC1414, 32'h010E261E, 32'h27FF1320, 32'h14FDEBCC, 
    /* (302, 0) */	    32'hC4C81515, 32'h010F2920, 32'h2AFF1422, 32'h16FDEAC8, 
    /* (303, 0) */	    32'hC0C41717, 32'h01102C22, 32'h2DFF1625, 32'h17FDE8C4, 
    /* (304, 0) */	    32'hBBC01818, 32'h01112F25, 32'h30FF1727, 32'h19FDE7C0, 
    /* (305, 0) */	    32'hB7BC1A1A, 32'h01123227, 32'h33FF1929, 32'h1AFCE5BC, 
    /* (306, 0) */	    32'hB3B81B1B, 32'h01133429, 32'h36FF1A2C, 32'h1CFCE3B8, 
    /* (307, 0) */	    32'hAFB41D1D, 32'h0114372B, 32'h39FF1C2E, 32'h1DFCE2B4, 
    /* (308, 0) */	    32'hAAB01F1F, 32'h01153A2E, 32'h3CFF1D31, 32'h1FFCE0B0, 
    /* (309, 0) */	    32'hA6AC2020, 32'h01163D30, 32'h3FFF1F33, 32'h20FCDFAC, 
    /* (310, 0) */	    32'hA2A82222, 32'h01174032, 32'h43FF2036, 32'h22FBDDA8, 
    /* (311, 0) */	    32'h9DA42323, 32'h01184335, 32'h46FF2238, 32'h23FBDBA4, 
    /* (312, 0) */	    32'h99A02525, 32'h011A4637, 32'h49FF233A, 32'h25FBDAA0, 
    /* (313, 0) */	    32'h959C2626, 32'h011B4939, 32'h4CFF243D, 32'h27FBD89C, 
    /* (314, 0) */	    32'h91982828, 32'h011C4C3B, 32'h4FFF263F, 32'h28FBD798, 
    /* (315, 0) */	    32'h8C942929, 32'h011D4F3E, 32'h52FF2742, 32'h2AFAD594, 
    /* (316, 0) */	    32'h88902B2B, 32'h011E5240, 32'h55FF2944, 32'h2BFAD390, 
    /* (317, 0) */	    32'h848C2C2C, 32'h011F5442, 32'h58FF2A47, 32'h2DFAD28C, 
    /* (318, 0) */	    32'h80892E2E, 32'h01205745, 32'h5BFF2C49, 32'h2EFAD088, 
    /* (319, 0) */	    32'h80852F2F, 32'h02215A47, 32'h5EFF2D4C, 32'h30FACF84, 
    /* (320, 0) */	    32'h84808013, 32'h7F018080, 32'h3E1C7C58, 32'h7F7FF769, 
    /* (321, 0) */	    32'h88848412, 32'h7C018484, 32'h3D1C7855, 32'h7C7CF866, 
    /* (322, 0) */	    32'h8C888812, 32'h78018888, 32'h3B1B7452, 32'h7878F863, 
    /* (323, 0) */	    32'h8F8C8C11, 32'h74018C8C, 32'h391A7050, 32'h7474F860, 
    /* (324, 0) */	    32'h93909011, 32'h70019090, 32'h37196C4D, 32'h7070F85C, 
    /* (325, 0) */	    32'h97949410, 32'h6C019494, 32'h3518684A, 32'h6C6CF959, 
    /* (326, 0) */	    32'h9B98980F, 32'h68019898, 32'h33176547, 32'h6868F956, 
    /* (327, 0) */	    32'h9F9C9C0F, 32'h64019C9C, 32'h31166145, 32'h6464F952, 
    /* (328, 0) */	    32'hA3A0A00E, 32'h6001A0A0, 32'h2F155D42, 32'h6060FA4F, 
    /* (329, 0) */	    32'hA7A4A40E, 32'h5C01A4A4, 32'h2D14593F, 32'h5C5CFA4C, 
    /* (330, 0) */	    32'hABA8A80D, 32'h5801A8A8, 32'h2B14553C, 32'h5858FA48, 
    /* (331, 0) */	    32'hAEACAC0C, 32'h5401ACAC, 32'h2913513A, 32'h5454FA45, 
    /* (332, 0) */	    32'hB2B0B00C, 32'h5001B0B0, 32'h27124D37, 32'h5050FB42, 
    /* (333, 0) */	    32'hB6B4B40B, 32'h4C01B4B4, 32'h25114934, 32'h4C4CFB3F, 
    /* (334, 0) */	    32'hBAB8B80B, 32'h4801B8B8, 32'h23104631, 32'h4848FB3B, 
    /* (335, 0) */	    32'hBEBCBC0A, 32'h4401BCBC, 32'h210F422F, 32'h4444FB38, 
    /* (336, 0) */	    32'hC2C0C009, 32'h4001C0C0, 32'h1F0E3E2C, 32'h4040FC35, 
    /* (337, 0) */	    32'hC6C4C409, 32'h3C01C4C4, 32'h1D0D3A29, 32'h3C3CFC31, 
    /* (338, 0) */	    32'hCAC8C808, 32'h3801C8C8, 32'h1B0C3626, 32'h3838FC2E, 
    /* (339, 0) */	    32'hCECCCC08, 32'h3400CCCC, 32'h190C3224, 32'h3434FD2B, 
    /* (340, 0) */	    32'hD1D0D007, 32'h3000D0D0, 32'h170B2E21, 32'h3030FD28, 
    /* (341, 0) */	    32'hD5D4D407, 32'h2C00D4D4, 32'h150A2B1E, 32'h2C2CFD24, 
    /* (342, 0) */	    32'hD9D8D806, 32'h2800D8D8, 32'h1409271B, 32'h2828FD21, 
    /* (343, 0) */	    32'hDDDCDC05, 32'h2400DCDC, 32'h12082319, 32'h2424FE1E, 
    /* (344, 0) */	    32'hE1E0E005, 32'h2000E0E0, 32'h10071F16, 32'h2020FE1A, 
    /* (345, 0) */	    32'hE5E4E404, 32'h1C00E4E4, 32'h0E061B13, 32'h1C1CFE17, 
    /* (346, 0) */	    32'hE9E8E804, 32'h1800E8E8, 32'h0C051710, 32'h1818FE14, 
    /* (347, 0) */	    32'hEDECEC03, 32'h1400ECEC, 32'h0A04130E, 32'h1414FF10, 
    /* (348, 0) */	    32'hF0F0F002, 32'h1000F0F0, 32'h08040F0B, 32'h1010FF0D, 
    /* (349, 0) */	    32'hF4F4F402, 32'h0C00F4F4, 32'h06030C08, 32'h0C0CFF0A, 
    /* (350, 0) */	    32'hF8F8F801, 32'h0800F8F8, 32'h04020805, 32'h0808FF07, 
    /* (351, 0) */	    32'hFCFCFC01, 32'h0400FCFC, 32'h02010403, 32'h04040003, 
    /* (352, 0) */	    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
    /* (353, 0) */	    32'h040404FF, 32'hFC000404, 32'hFEFFFCFD, 32'hFCFC00FD, 
    /* (354, 0) */	    32'h080808FF, 32'hF8000808, 32'hFCFEF8FB, 32'hF8F801F9, 
    /* (355, 0) */	    32'h0C0C0CFE, 32'hF4000C0C, 32'hFAFDF4F8, 32'hF4F401F6, 
    /* (356, 0) */	    32'h101010FE, 32'hF0001010, 32'hF8FCF1F5, 32'hF0F001F3, 
    /* (357, 0) */	    32'h131414FD, 32'hEC001414, 32'hF6FCEDF2, 32'hECEC01F0, 
    /* (358, 0) */	    32'h171818FC, 32'hE8001818, 32'hF4FBE9F0, 32'hE8E802EC, 
    /* (359, 0) */	    32'h1B1C1CFC, 32'hE4001C1C, 32'hF2FAE5ED, 32'hE4E402E9, 
    /* (360, 0) */	    32'h1F2020FB, 32'hE0002020, 32'hF0F9E1EA, 32'hE0E002E6, 
    /* (361, 0) */	    32'h232424FB, 32'hDC002424, 32'hEEF8DDE7, 32'hDCDC02E2, 
    /* (362, 0) */	    32'h272828FA, 32'hD8002828, 32'hECF7D9E5, 32'hD8D803DF, 
    /* (363, 0) */	    32'h2B2C2CF9, 32'hD4002C2C, 32'hEBF6D5E2, 32'hD4D403DC, 
    /* (364, 0) */	    32'h2F3030F9, 32'hD0003030, 32'hE9F5D2DF, 32'hD0D003D8, 
    /* (365, 0) */	    32'h323434F8, 32'hCC003434, 32'hE7F4CEDC, 32'hCCCC03D5, 
    /* (366, 0) */	    32'h363838F8, 32'hC8FF3838, 32'hE5F4CADA, 32'hC8C804D2, 
    /* (367, 0) */	    32'h3A3C3CF7, 32'hC4FF3C3C, 32'hE3F3C6D7, 32'hC4C404CF, 
    /* (368, 0) */	    32'h3E4040F7, 32'hC0FF4040, 32'hE1F2C2D4, 32'hC0C004CB, 
    /* (369, 0) */	    32'h424444F6, 32'hBCFF4444, 32'hDFF1BED1, 32'hBCBC05C8, 
    /* (370, 0) */	    32'h464848F5, 32'hB8FF4848, 32'hDDF0BACF, 32'hB8B805C5, 
    /* (371, 0) */	    32'h4A4C4CF5, 32'hB4FF4C4C, 32'hDBEFB7CC, 32'hB4B405C1, 
    /* (372, 0) */	    32'h4E5050F4, 32'hB0FF5050, 32'hD9EEB3C9, 32'hB0B005BE, 
    /* (373, 0) */	    32'h525454F4, 32'hACFF5454, 32'hD7EDAFC6, 32'hACAC06BB, 
    /* (374, 0) */	    32'h555858F3, 32'hA8FF5858, 32'hD5ECABC4, 32'hA8A806B8, 
    /* (375, 0) */	    32'h595C5CF2, 32'hA4FF5C5C, 32'hD3ECA7C1, 32'hA4A406B4, 
    /* (376, 0) */	    32'h5D6060F2, 32'hA0FF6060, 32'hD1EBA3BE, 32'hA0A006B1, 
    /* (377, 0) */	    32'h616464F1, 32'h9CFF6464, 32'hCFEA9FBB, 32'h9C9C07AE, 
    /* (378, 0) */	    32'h656868F1, 32'h98FF6868, 32'hCDE99BB9, 32'h989807AA, 
    /* (379, 0) */	    32'h696C6CF0, 32'h94FF6C6C, 32'hCBE898B6, 32'h949407A7, 
    /* (380, 0) */	    32'h6D7070EF, 32'h90FF7070, 32'hC9E794B3, 32'h909008A4, 
    /* (381, 0) */	    32'h717474EF, 32'h8CFF7474, 32'hC7E690B0, 32'h8C8C08A0, 
    /* (382, 0) */	    32'h747878EE, 32'h88FF7878, 32'hC5E58CAE, 32'h8888089D, 
    /* (383, 0) */	    32'h787C7CEE, 32'h84FF7C7C, 32'hC3E488AB, 32'h8484089A, 
    /* (384, 0) */	    32'h25C10373, 32'hE8DBF2E7, 32'hB710ED1B, 32'hF5DE2103, 
    /* (385, 0) */	    32'h24C30370, 32'hE9DCF2E8, 32'hB910EE1A, 32'hF5DF2003, 
    /* (386, 0) */	    32'h23C5036C, 32'hEADDF3E9, 32'hBC0FEE19, 32'hF6E01F03, 
    /* (387, 0) */	    32'h22C70369, 32'hEBDEF3E9, 32'hBE0FEF18, 32'hF6E11E03, 
    /* (388, 0) */	    32'h21C90365, 32'hEBE0F4EA, 32'hC00EF017, 32'hF6E21D03, 
    /* (389, 0) */	    32'h20CB0361, 32'hECE1F4EB, 32'hC30EF016, 32'hF7E31C03, 
    /* (390, 0) */	    32'h1ECD035E, 32'hEDE2F4EC, 32'hC50DF116, 32'hF7E41B02, 
    /* (391, 0) */	    32'h1DCF035A, 32'hEEE3F5ED, 32'hC70DF115, 32'hF7E51A02, 
    /* (392, 0) */	    32'h1CD10257, 32'hEEE4F5ED, 32'hC90CF214, 32'hF8E61902, 
    /* (393, 0) */	    32'h1BD30253, 32'hEFE5F6EE, 32'hCC0CF313, 32'hF8E71802, 
    /* (394, 0) */	    32'h1AD5024F, 32'hF0E7F6EF, 32'hCE0BF312, 32'hF8E91702, 
    /* (395, 0) */	    32'h19D7024C, 32'hF1E8F7F0, 32'hD00BF411, 32'hF9EA1602, 
    /* (396, 0) */	    32'h17D90248, 32'hF1E9F7F0, 32'hD20AF411, 32'hF9EB1502, 
    /* (397, 0) */	    32'h16DB0244, 32'hF2EAF8F1, 32'hD50AF510, 32'hF9EC1402, 
    /* (398, 0) */	    32'h15DC0241, 32'hF3EBF8F2, 32'hD709F50F, 32'hFAED1302, 
    /* (399, 0) */	    32'h14DE023D, 32'hF3ECF8F3, 32'hD909F60E, 32'hFAEE1202, 
    /* (400, 0) */	    32'h13E0023A, 32'hF4EDF9F4, 32'hDC08F70D, 32'hFBEF1101, 
    /* (401, 0) */	    32'h12E20236, 32'hF5EFF9F4, 32'hDE08F70C, 32'hFBF01001, 
    /* (402, 0) */	    32'h10E40132, 32'hF6F0FAF5, 32'hE007F80C, 32'hFBF10E01, 
    /* (403, 0) */	    32'h0FE6012F, 32'hF6F1FAF6, 32'hE207F80B, 32'hFCF20D01, 
    /* (404, 0) */	    32'h0EE8012B, 32'hF7F2FBF7, 32'hE506F90A, 32'hFCF30C01, 
    /* (405, 0) */	    32'h0DEA0128, 32'hF8F3FBF7, 32'hE706FA09, 32'hFCF40B01, 
    /* (406, 0) */	    32'h0CEC0124, 32'hF9F4FCF8, 32'hE905FA08, 32'hFDF50A01, 
    /* (407, 0) */	    32'h0BEE0120, 32'hF9F6FCF9, 32'hEC05FB07, 32'hFDF60901, 
    /* (408, 0) */	    32'h09F0011D, 32'hFAF7FCFA, 32'hEE04FB07, 32'hFDF70801, 
    /* (409, 0) */	    32'h08F20119, 32'hFBF8FDFB, 32'hF004FC06, 32'hFEF90701, 
    /* (410, 0) */	    32'h07F40116, 32'hFCF9FDFB, 32'hF203FC05, 32'hFEFA0601, 
    /* (411, 0) */	    32'h06F60112, 32'hFCFAFEFC, 32'hF503FD04, 32'hFEFB0500, 
    /* (412, 0) */	    32'h05F8000E, 32'hFDFBFEFD, 32'hF702FE03, 32'hFFFC0400, 
    /* (413, 0) */	    32'h04FA000B, 32'hFEFDFFFE, 32'hF902FE02, 32'hFFFD0300, 
    /* (414, 0) */	    32'h02FC0007, 32'hFFFEFFFE, 32'hFB01FF02, 32'hFFFE0200, 
    /* (415, 0) */	    32'h01FE0004, 32'hFFFF00FF, 32'hFE01FF01, 32'h00FF0100, 
    /* (416, 0) */	    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
    /* (417, 0) */	    32'hFF0200FC, 32'h01010001, 32'h02FF01FF, 32'h0001FF00, 
    /* (418, 0) */	    32'hFE0400F9, 32'h01020102, 32'h05FF01FE, 32'h0102FE00, 
    /* (419, 0) */	    32'hFC0600F5, 32'h02030102, 32'h07FE02FE, 32'h0103FD00, 
    /* (420, 0) */	    32'hFB0800F2, 32'h03050203, 32'h09FE02FD, 32'h0104FC00, 
    /* (421, 0) */	    32'hFA0AFFEE, 32'h04060204, 32'h0BFD03FC, 32'h0205FB00, 
    /* (422, 0) */	    32'hF90CFFEA, 32'h04070305, 32'h0EFD04FB, 32'h0206FAFF, 
    /* (423, 0) */	    32'hF80EFFE7, 32'h05080305, 32'h10FC04FA, 32'h0207F9FF, 
    /* (424, 0) */	    32'hF710FFE3, 32'h06090406, 32'h12FC05F9, 32'h0309F8FF, 
    /* (425, 0) */	    32'hF512FFE0, 32'h070A0407, 32'h14FB05F9, 32'h030AF7FF, 
    /* (426, 0) */	    32'hF414FFDC, 32'h070C0408, 32'h17FB06F8, 32'h030BF6FF, 
    /* (427, 0) */	    32'hF316FFD8, 32'h080D0509, 32'h19FA06F7, 32'h040CF5FF, 
    /* (428, 0) */	    32'hF218FFD5, 32'h090E0509, 32'h1BFA07F6, 32'h040DF4FF, 
    /* (429, 0) */	    32'hF11AFFD1, 32'h0A0F060A, 32'h1EF908F5, 32'h040EF3FF, 
    /* (430, 0) */	    32'hF01CFFCE, 32'h0A10060B, 32'h20F908F4, 32'h050FF2FF, 
    /* (431, 0) */	    32'hEE1EFECA, 32'h0B11070C, 32'h22F809F4, 32'h0510F0FF, 
    /* (432, 0) */	    32'hED20FEC6, 32'h0C13070C, 32'h24F809F3, 32'h0511EFFF, 
    /* (433, 0) */	    32'hEC22FEC3, 32'h0D14080D, 32'h27F70AF2, 32'h0612EEFE, 
    /* (434, 0) */	    32'hEB24FEBF, 32'h0D15080E, 32'h29F70BF1, 32'h0613EDFE, 
    /* (435, 0) */	    32'hEA25FEBC, 32'h0E16080F, 32'h2BF60BF0, 32'h0714ECFE, 
    /* (436, 0) */	    32'hE927FEB8, 32'h0F170910, 32'h2EF60CEF, 32'h0715EBFE, 
    /* (437, 0) */	    32'hE729FEB4, 32'h0F180910, 32'h30F50CEF, 32'h0716EAFE, 
    /* (438, 0) */	    32'hE62BFEB1, 32'h10190A11, 32'h32F50DEE, 32'h0817E9FE, 
    /* (439, 0) */	    32'hE52DFEAD, 32'h111B0A12, 32'h34F40DED, 32'h0819E8FE, 
    /* (440, 0) */	    32'hE42FFEA9, 32'h121C0B13, 32'h37F40EEC, 32'h081AE7FE, 
    /* (441, 0) */	    32'hE331FDA6, 32'h121D0B13, 32'h39F30FEB, 32'h091BE6FE, 
    /* (442, 0) */	    32'hE233FDA2, 32'h131E0C14, 32'h3BF30FEA, 32'h091CE5FE, 
    /* (443, 0) */	    32'hE035FD9F, 32'h141F0C15, 32'h3DF210EA, 32'h091DE4FD, 
    /* (444, 0) */	    32'hDF37FD9B, 32'h15200C16, 32'h40F210E9, 32'h0A1EE3FD, 
    /* (445, 0) */	    32'hDE39FD97, 32'h15220D17, 32'h42F111E8, 32'h0A1FE2FD, 
    /* (446, 0) */	    32'hDD3BFD94, 32'h16230D17, 32'h44F112E7, 32'h0A20E1FD, 
    /* (447, 0) */	    32'hDC3DFD90, 32'h17240E18, 32'h47F012E6, 32'h0B21E0FD, 
    /* (448, 0) */	    32'hDC7F4280, 32'h2970505E, 32'h7F7F7F80, 32'h317F8080, 
    /* (449, 0) */	    32'hDD7C4080, 32'h276D4D5C, 32'h7C7B7C84, 32'h307B8484, 
    /* (450, 0) */	    32'hDE783E84, 32'h26694B59, 32'h78777888, 32'h2E778888, 
    /* (451, 0) */	    32'hDF743B88, 32'h25664856, 32'h7473748C, 32'h2D748C8C, 
    /* (452, 0) */	    32'hE070398D, 32'h24624653, 32'h70707090, 32'h2B709090, 
    /* (453, 0) */	    32'hE16C3791, 32'h225F4350, 32'h6C6C6C94, 32'h296C9494, 
    /* (454, 0) */	    32'hE3683595, 32'h215B414D, 32'h68686898, 32'h28689898, 
    /* (455, 0) */	    32'hE4643399, 32'h20583E4A, 32'h6464649C, 32'h26649C9C, 
    /* (456, 0) */	    32'hE560319D, 32'h1E543C47, 32'h606060A0, 32'h2560A0A0, 
    /* (457, 0) */	    32'hE65C2FA1, 32'h1D513944, 32'h5C5C5CA4, 32'h235CA4A4, 
    /* (458, 0) */	    32'hE7582DA5, 32'h1C4D3741, 32'h585858A8, 32'h2258A8A8, 
    /* (459, 0) */	    32'hE8542BA9, 32'h1B4A343E, 32'h545454AC, 32'h2054ACAC, 
    /* (460, 0) */	    32'hE95029AE, 32'h1946323B, 32'h505050B0, 32'h1F50B0B0, 
    /* (461, 0) */	    32'hEB4C27B2, 32'h18432F38, 32'h4C4C4CB4, 32'h1D4CB4B4, 
    /* (462, 0) */	    32'hEC4825B6, 32'h173F2D35, 32'h484848B8, 32'h1C48B8B8, 
    /* (463, 0) */	    32'hED4423BA, 32'h163C2A32, 32'h444444BC, 32'h1A44BCBC, 
    /* (464, 0) */	    32'hEE4021BE, 32'h1438282F, 32'h404040C0, 32'h1940C0C0, 
    /* (465, 0) */	    32'hEF3C1FC2, 32'h1335252C, 32'h3C3C3CC4, 32'h173CC4C4, 
    /* (466, 0) */	    32'hF0381DC6, 32'h12312329, 32'h383838C8, 32'h1638C8C8, 
    /* (467, 0) */	    32'hF1341BCA, 32'h112E2026, 32'h343434CC, 32'h1434CCCC, 
    /* (468, 0) */	    32'hF23019CF, 32'h0F2A1E23, 32'h303030D0, 32'h1230D0D0, 
    /* (469, 0) */	    32'hF42C17D3, 32'h0E271B20, 32'h2C2C2CD4, 32'h112CD4D4, 
    /* (470, 0) */	    32'hF52815D7, 32'h0D23191E, 32'h282828D8, 32'h0F28D8D8, 
    /* (471, 0) */	    32'hF62412DB, 32'h0B20161B, 32'h242424DC, 32'h0E24DCDC, 
    /* (472, 0) */	    32'hF72010DF, 32'h0A1C1418, 32'h202020E0, 32'h0C20E0E0, 
    /* (473, 0) */	    32'hF81C0EE3, 32'h09191115, 32'h1C1C1CE4, 32'h0B1CE4E4, 
    /* (474, 0) */	    32'hF9180CE7, 32'h08150F12, 32'h181818E8, 32'h0918E8E8, 
    /* (475, 0) */	    32'hFA140AEB, 32'h06120C0F, 32'h141414EC, 32'h0814ECEC, 
    /* (476, 0) */	    32'hFB1008F0, 32'h050E0A0C, 32'h101010F0, 32'h0610F0F0, 
    /* (477, 0) */	    32'hFD0C06F4, 32'h040B0709, 32'h0C0C0CF4, 32'h050CF4F4, 
    /* (478, 0) */	    32'hFE0804F8, 32'h03070506, 32'h080808F8, 32'h0308F8F8, 
    /* (479, 0) */	    32'hFF0402FC, 32'h01040203, 32'h040404FC, 32'h0204FCFC, 
    /* (480, 0) */	    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
    /* (481, 0) */	    32'h01FCFE04, 32'hFFFCFEFD, 32'hFCFCFC04, 32'hFEFC0404, 
    /* (482, 0) */	    32'h02F8FC08, 32'hFDF9FBFA, 32'hF8F8F808, 32'hFDF80808, 
    /* (483, 0) */	    32'h03F4FA0C, 32'hFCF5F9F7, 32'hF4F4F40C, 32'hFBF40C0C, 
    /* (484, 0) */	    32'h05F0F810, 32'hFBF2F6F4, 32'hF0F0F010, 32'hFAF01010, 
    /* (485, 0) */	    32'h06ECF615, 32'hFAEEF4F1, 32'hECECEC14, 32'hF8EC1414, 
    /* (486, 0) */	    32'h07E8F419, 32'hF8EBF1EE, 32'hE8E8E818, 32'hF7E81818, 
    /* (487, 0) */	    32'h08E4F21D, 32'hF7E7EFEB, 32'hE4E4E41C, 32'hF5E41C1C, 
    /* (488, 0) */	    32'h09E0F021, 32'hF6E4ECE8, 32'hE0E0E020, 32'hF4E02020, 
    /* (489, 0) */	    32'h0ADCEE25, 32'hF5E0EAE5, 32'hDCDCDC24, 32'hF2DC2424, 
    /* (490, 0) */	    32'h0BD8EB29, 32'hF3DDE7E2, 32'hD8D8D828, 32'hF1D82828, 
    /* (491, 0) */	    32'h0CD4E92D, 32'hF2D9E5E0, 32'hD4D4D42C, 32'hEFD42C2C, 
    /* (492, 0) */	    32'h0ED0E731, 32'hF1D6E2DD, 32'hD0D0D030, 32'hEED03030, 
    /* (493, 0) */	    32'h0FCCE536, 32'hEFD2E0DA, 32'hCCCCCC34, 32'hECCC3434, 
    /* (494, 0) */	    32'h10C8E33A, 32'hEECFDDD7, 32'hC8C8C838, 32'hEAC83838, 
    /* (495, 0) */	    32'h11C4E13E, 32'hEDCBDBD4, 32'hC4C4C43C, 32'hE9C43C3C, 
    /* (496, 0) */	    32'h12C0DF42, 32'hECC8D8D1, 32'hC0C0C040, 32'hE7C04040, 
    /* (497, 0) */	    32'h13BCDD46, 32'hEAC4D6CE, 32'hBCBCBC44, 32'hE6BC4444, 
    /* (498, 0) */	    32'h14B8DB4A, 32'hE9C1D3CB, 32'hB8B8B848, 32'hE4B84848, 
    /* (499, 0) */	    32'h15B4D94E, 32'hE8BDD1C8, 32'hB4B4B44C, 32'hE3B44C4C, 
    /* (500, 0) */	    32'h17B0D752, 32'hE7BACEC5, 32'hB0B0B050, 32'hE1B05050, 
    /* (501, 0) */	    32'h18ACD557, 32'hE5B6CCC2, 32'hACACAC54, 32'hE0AC5454, 
    /* (502, 0) */	    32'h19A8D35B, 32'hE4B3C9BF, 32'hA8A8A858, 32'hDEA85858, 
    /* (503, 0) */	    32'h1AA4D15F, 32'hE3AFC7BC, 32'hA4A4A45C, 32'hDDA45C5C, 
    /* (504, 0) */	    32'h1BA0CF63, 32'hE2ACC4B9, 32'hA0A0A060, 32'hDBA06060, 
    /* (505, 0) */	    32'h1C9CCD67, 32'hE0A8C2B6, 32'h9C9C9C64, 32'hDA9C6464, 
    /* (506, 0) */	    32'h1D98CB6B, 32'hDFA5BFB3, 32'h98989868, 32'hD8986868, 
    /* (507, 0) */	    32'h1F94C96F, 32'hDEA1BDB0, 32'h9494946C, 32'hD7946C6C, 
    /* (508, 0) */	    32'h2090C773, 32'hDC9EBAAD, 32'h90909070, 32'hD5907070, 
    /* (509, 0) */	    32'h218CC578, 32'hDB9AB8AA, 32'h8C8D8C74, 32'hD38C7474, 
    /* (510, 0) */	    32'h2288C27C, 32'hDA97B5A7, 32'h88898878, 32'hD2897878, 
    /* (511, 0) */	    32'h2384C07F, 32'hD993B3A4, 32'h8485847C, 32'hD0857C7C, 
    /* (512, 0) */	    32'h7F354F7F, 32'h4E7F7F7F, 32'h177BC57F, 32'h7C7F2E7F, 
    /* (513, 0) */	    32'h7F344D7F, 32'h4B7F7F7F, 32'h1777C67F, 32'h797F2C7F, 
    /* (514, 0) */	    32'h7F324B7F, 32'h497F7F7F, 32'h1673C87F, 32'h757F2B7F, 
    /* (515, 0) */	    32'h7F30487F, 32'h467C7F7F, 32'h156FCA7C, 32'h717F2A7D, 
    /* (516, 0) */	    32'h7F2F467F, 32'h44787F7F, 32'h156CCC78, 32'h6D7F2879, 
    /* (517, 0) */	    32'h7F2D437F, 32'h42737F7F, 32'h1468CE74, 32'h697F2775, 
    /* (518, 0) */	    32'h7F2B417F, 32'h3F6F7F7F, 32'h1364D06F, 32'h657F2570, 
    /* (519, 0) */	    32'h7F2A3E7F, 32'h3D6B7F7F, 32'h1260D26B, 32'h617F246C, 
    /* (520, 0) */	    32'h7F283C7F, 32'h3A677F7F, 32'h125CD367, 32'h5D7D2268, 
    /* (521, 0) */	    32'h7F26397F, 32'h38627F7F, 32'h1158D563, 32'h59782163, 
    /* (522, 0) */	    32'h7F25377F, 32'h355E7F7D, 32'h1055D75E, 32'h5673205F, 
    /* (523, 0) */	    32'h7F23347F, 32'h335A7F77, 32'h0F51D95A, 32'h526D1E5B, 
    /* (524, 0) */	    32'h7F21327F, 32'h31557F71, 32'h0F4DDB56, 32'h4E681D56, 
    /* (525, 0) */	    32'h7F202F7F, 32'h2E517F6C, 32'h0E49DD51, 32'h4A631B52, 
    /* (526, 0) */	    32'h7F1E2D7F, 32'h2C4D7C66, 32'h0D45DF4D, 32'h465E1A4E, 
    /* (527, 0) */	    32'h781C2A7F, 32'h29497560, 32'h0C41E049, 32'h42591849, 
    /* (528, 0) */	    32'h711B287F, 32'h27446E5B, 32'h0C3DE245, 32'h3E531745, 
    /* (529, 0) */	    32'h6A19257F, 32'h24406755, 32'h0B3AE440, 32'h3A4E1541, 
    /* (530, 0) */	    32'h6317237C, 32'h223C604F, 32'h0A36E63C, 32'h3649143C, 
    /* (531, 0) */	    32'h5C162073, 32'h2038594A, 32'h0A32E838, 32'h33441338, 
    /* (532, 0) */	    32'h55141E6A, 32'h1D335244, 32'h092EEA33, 32'h2F3E1134, 
    /* (533, 0) */	    32'h4E121B61, 32'h1B2F4C3E, 32'h082AEC2F, 32'h2B39102F, 
    /* (534, 0) */	    32'h47111958, 32'h182B4539, 32'h0726ED2B, 32'h27340E2B, 
    /* (535, 0) */	    32'h3F0F164F, 32'h16263E33, 32'h0723EF27, 32'h232F0D27, 
    /* (536, 0) */	    32'h380D1447, 32'h1322372D, 32'h061FF122, 32'h1F2A0B23, 
    /* (537, 0) */	    32'h310C113E, 32'h111E3028, 32'h051BF31E, 32'h1B240A1E, 
    /* (538, 0) */	    32'h2A0A0F35, 32'h0F1A2922, 32'h0417F51A, 32'h171F091A, 
    /* (539, 0) */	    32'h23080C2C, 32'h0C15221C, 32'h0413F715, 32'h131A0716, 
    /* (540, 0) */	    32'h1C070A23, 32'h0A111B17, 32'h030FF911, 32'h10150611, 
    /* (541, 0) */	    32'h1505071A, 32'h070D1511, 32'h020CFA0D, 32'h0C10040D, 
    /* (542, 0) */	    32'h0E030512, 32'h05090E0B, 32'h0108FC09, 32'h080A0309, 
    /* (543, 0) */	    32'h07020209, 32'h02040706, 32'h0104FE04, 32'h04050104, 
    /* (544, 0) */	    32'h00000000, 32'h00000000, 32'h00000000, 32'h00000000, 
    /* (545, 0) */	    32'hF9FEFEF7, 32'hFEFCF9FA, 32'hFFFC02FC, 32'hFCFBFFFC, 
    /* (546, 0) */	    32'hF2FDFBEE, 32'hFBF7F2F5, 32'hFFF804F7, 32'hF8F6FDF7, 
    /* (547, 0) */	    32'hEBFBF9E6, 32'hF9F3EBEF, 32'hFEF406F3, 32'hF4F0FCF3, 
    /* (548, 0) */	    32'hE4F9F6DD, 32'hF6EFE5E9, 32'hFDF107EF, 32'hF0EBFAEF, 
    /* (549, 0) */	    32'hDDF8F4D4, 32'hF4EBDEE4, 32'hFCED09EB, 32'hEDE6F9EA, 
    /* (550, 0) */	    32'hD6F6F1CB, 32'hF1E6D7DE, 32'hFCE90BE6, 32'hE9E1F7E6, 
    /* (551, 0) */	    32'hCFF4EFC2, 32'hEFE2D0D8, 32'hFBE50DE2, 32'hE5DCF6E2, 
    /* (552, 0) */	    32'hC8F3ECB9, 32'hEDDEC9D3, 32'hFAE10FDE, 32'hE1D6F5DD, 
    /* (553, 0) */	    32'hC1F1EAB1, 32'hEADAC2CD, 32'hF9DD11D9, 32'hDDD1F3D9, 
    /* (554, 0) */	    32'hB9EFE7A8, 32'hE8D5BBC7, 32'hF9DA13D5, 32'hD9CCF2D5, 
    /* (555, 0) */	    32'hB2EEE59F, 32'hE5D1B4C2, 32'hF8D614D1, 32'hD5C7F0D1, 
    /* (556, 0) */	    32'hABECE296, 32'hE3CDAEBC, 32'hF7D216CD, 32'hD1C2EFCC, 
    /* (557, 0) */	    32'hA4EAE08D, 32'hE0C8A7B6, 32'hF6CE18C8, 32'hCDBCEDC8, 
    /* (558, 0) */	    32'h9DE9DD84, 32'hDEC4A0B1, 32'hF6CA1AC4, 32'hCAB7ECC4, 
    /* (559, 0) */	    32'h96E7DB80, 32'hDCC099AB, 32'hF5C61CC0, 32'hC6B2EBBF, 
    /* (560, 0) */	    32'h8FE5D880, 32'hD9BC92A5, 32'hF4C31EBB, 32'hC2ADE9BB, 
    /* (561, 0) */	    32'h88E4D680, 32'hD7B78BA0, 32'hF4BF20B7, 32'hBEA7E8B7, 
    /* (562, 0) */	    32'h81E2D380, 32'hD4B3849A, 32'hF3BB21B3, 32'hBAA2E6B2, 
    /* (563, 0) */	    32'h80E0D180, 32'hD2AF8094, 32'hF2B723AF, 32'hB69DE5AE, 
    /* (564, 0) */	    32'h80DFCE80, 32'hCFAB808F, 32'hF1B325AA, 32'hB298E3AA, 
    /* (565, 0) */	    32'h80DDCC80, 32'hCDA68089, 32'hF1AF27A6, 32'hAE93E2A5, 
    /* (566, 0) */	    32'h80DBC980, 32'hCBA28083, 32'hF0AB29A2, 32'hAA8DE0A1, 
    /* (567, 0) */	    32'h80DAC780, 32'hC89E8080, 32'hEFA82B9D, 32'hA788DF9D, 
    /* (568, 0) */	    32'h80D8C480, 32'hC6998080, 32'hEEA42D99, 32'hA383DE98, 
    /* (569, 0) */	    32'h80D6C280, 32'hC3958080, 32'hEEA02E95, 32'h9F80DC94, 
    /* (570, 0) */	    32'h80D5BF80, 32'hC1918080, 32'hED9C3091, 32'h9B80DB90, 
    /* (571, 0) */	    32'h80D3BD80, 32'hBE8D8080, 32'hEC98328C, 32'h9780D98B, 
    /* (572, 0) */	    32'h80D1BA80, 32'hBC888080, 32'hEB943488, 32'h9380D887, 
    /* (573, 0) */	    32'h80D0B880, 32'hBA848080, 32'hEB913684, 32'h8F80D683, 
    /* (574, 0) */	    32'h80CEB580, 32'hB7808080, 32'hEA8D3880, 32'h8B80D580, 
    /* (575, 0) */	    32'h80CCB380, 32'hB5808080, 32'hE9893A80, 32'h8780D480
};

    // 写入数据
    always_latch begin
        if (en_write) begin
            lut_mem[base * 4 + 0] = wdata[0];
            lut_mem[base * 4 + 1] = wdata[1];
            lut_mem[base * 4 + 2] = wdata[2];
            lut_mem[base * 4 + 3] = wdata[3];
        end else begin
            ;
        end
    end

    // 读取数据
    always_latch begin
        if (en_read) begin
            rdata[0] = lut_mem[base * 4 + 0];
            rdata[1] = lut_mem[base * 4 + 1];
            rdata[2] = lut_mem[base * 4 + 2];
            rdata[3] = lut_mem[base * 4 + 3];
        end else begin
            ;
        end
    end

endmodule
